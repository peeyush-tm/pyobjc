/*
 * WARNING: This is a generated file, do not change
 */

#include <Python.h>
#include <objc/objc.h>
#include <objc/objc-runtime.h>
#include <Foundation/NSException.h>
#define PYOBJC_METHOD_STUB_IMPL
#include "pyobjc-api.h"
static struct pyobjc_api* ObjC_API;
typedef int (*superfunc)();
/* signature: #12@4:8@12@16 */
static Class 
meth_imp_0(id self, SEL sel, id arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	Class objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("#", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_0(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	Class objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (Class)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("#", &objc_retval);
	return v;
}


/* signature: #4@4:8 */
static Class 
meth_imp_1(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	Class objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("#", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_1(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	Class objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (Class)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("#", &objc_retval);
	return v;
}


/* signature: #8@4:8@12 */
static Class 
meth_imp_2(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	Class objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("#", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_2(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	Class objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (Class)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("#", &objc_retval);
	return v;
}


/* signature: #8@4:8I12 */
static Class 
meth_imp_3(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	Class objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("#", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_3(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	Class objc_retval;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (Class)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("#", &objc_retval);
	return v;
}


/* signature: *12@4:8@12^I16 */
static char* 
meth_imp_4(id self, SEL sel, id arg_2, unsigned int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char* objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("*", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_4(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_retval;
	id objc_arg2;
	unsigned int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char*)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("*", &objc_retval);
	return v;
}


/* signature: *4@4:8 */
static char* 
meth_imp_5(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char* objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("*", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_5(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (char*)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("*", &objc_retval);
	return v;
}


/* signature: *8@4:8r*12 */
static char* 
meth_imp_6(id self, SEL sel, char* arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char* objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("*", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_6(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_retval;
	char* objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char*)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("*", &objc_retval);
	return v;
}


/* signature: :4@4:8 */
static SEL 
meth_imp_7(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	SEL objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC(":", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_7(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	SEL objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (SEL)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython(":", &objc_retval);
	return v;
}


/* signature: :8@4:8@12 */
static SEL 
meth_imp_8(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	SEL objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC(":", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_8(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	SEL objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (SEL)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython(":", &objc_retval);
	return v;
}


/* signature: @10@4:8S12S16 */
static id 
meth_imp_9(id self, SEL sel, unsigned short arg_2, unsigned short arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_9(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned short objc_arg2;
	unsigned short objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @120@4:8{_CGSEventRecord=SSII{CGPoint=ff}{CGPoint=ff}QI^v^v(?={?=CCsiCcCCss(?={_CGSTabletPointData=iiiSS{?=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})[4i]}{?=CCsiCcCCss(?={_CGSTabletPointData=iiiSS{?=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})[4i]}{?=ssSSSsssI[11i]}{?=ssii[13i]}{?=SSIIi[12i]}{?=ssssi[13i]}{?=iiiSS{?=ss}SsSsss[8i]}{?=SSSSSSIQICCs[8i]}{?=ss(?=[15f][15i][30s][60c])})}16 */
struct CGPoint {
	float field_0;
	float field_1;
};
struct pyobjcanonymous0 {
	short field_0;
	short field_1;
};
struct _CGSTabletPointData {
	int field_0;
	int field_1;
	int field_2;
	unsigned short field_3;
	unsigned short field_4;
	struct pyobjcanonymous0 field_5;
	unsigned short field_6;
	short field_7;
	unsigned short field_8;
	short field_9;
	short field_10;
	short field_11;
};
struct _CGSTabletProximityData {
	unsigned short field_0;
	unsigned short field_1;
	unsigned short field_2;
	unsigned short field_3;
	unsigned short field_4;
	unsigned short field_5;
	unsigned int field_6;
	unsigned long long field_7;
	unsigned int field_8;
	unsigned char field_9;
	unsigned char field_10;
	short field_11;
};
union pyobjcanonymous1 {	struct _CGSTabletPointData field_0;	struct _CGSTabletProximityData field_1;};
struct _CGSEventRecord {
	unsigned short field_0;
	unsigned short field_1;
	unsigned int field_2;
	unsigned int field_3;
	struct CGPoint field_4;
	struct CGPoint field_5;
	unsigned long long field_6;
	unsigned int field_7;
	void  *field_8;
	void  *field_9;
	union pyobjcanonymous1 field_10;
};

static id 
meth_imp_10(id self, SEL sel, struct _CGSEventRecord arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_CGSEventRecord=SSII{CGPoint=ff}{CGPoint=ff}QI^v^v(pyobjcanonymous1={_CGSTabletPointData=iiiSS{pyobjcanonymous0=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_10(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _CGSEventRecord objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_CGSEventRecord=SSII{CGPoint=ff}{CGPoint=ff}QI^v^v(pyobjcanonymous1={_CGSTabletPointData=iiiSS{pyobjcanonymous0=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @124@4:8{_CGSEventRecord=SSII{CGPoint=ff}{CGPoint=ff}QI^v^v(?={?=CCsiCcCCss(?={_CGSTabletPointData=iiiSS{?=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})[4i]}{?=CCsiCcCCss(?={_CGSTabletPointData=iiiSS{?=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})[4i]}{?=ssSSSsssI[11i]}{?=ssii[13i]}{?=SSIIi[12i]}{?=ssssi[13i]}{?=iiiSS{?=ss}SsSsss[8i]}{?=SSSSSSIQICCs[8i]}{?=ss(?=[15f][15i][30s][60c])})}16^v128 */
static id 
meth_imp_11(id self, SEL sel, struct _CGSEventRecord arg_2, void  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_CGSEventRecord=SSII{CGPoint=ff}{CGPoint=ff}QI^v^v(pyobjcanonymous1={_CGSTabletPointData=iiiSS{pyobjcanonymous0=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_11(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _CGSEventRecord objc_arg2;
	void  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_CGSEventRecord=SSII{CGPoint=ff}{CGPoint=ff}QI^v^v(pyobjcanonymous1={_CGSTabletPointData=iiiSS{pyobjcanonymous0=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8*12I16 */
static id 
meth_imp_12(id self, SEL sel, char* arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_12(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8*12i16 */
static id 
meth_imp_13(id self, SEL sel, char* arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_13(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8*16 */
static id 
meth_imp_14(id self, SEL sel, char* arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_14(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8:12@16 */
static id 
meth_imp_15(id self, SEL sel, SEL arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_15(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	SEL objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8:12^:16 */
static id 
meth_imp_16(id self, SEL sel, SEL arg_2, SEL  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^:", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_16(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	SEL objc_arg2;
	SEL  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^:", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8:12^v16 */
static id 
meth_imp_17(id self, SEL sel, SEL arg_2, void  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_17(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	SEL objc_arg2;
	void  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8@12#16 */
static id 
meth_imp_18(id self, SEL sel, id arg_2, Class arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_18(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	Class objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8@12*16 */
static id 
meth_imp_19(id self, SEL sel, id arg_2, char* arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_19(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	char* objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8@12@16 */
static id 
meth_imp_20(id self, SEL sel, id arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_20(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8@12I16 */
static id 
meth_imp_21(id self, SEL sel, id arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_21(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8@12^{?=^SI^SI^SI}16 */
static id 
meth_imp_22(id self, SEL sel, id arg_2, struct pyobjcanonymous0  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_22(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct pyobjcanonymous0  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8@12^{_NSZone=}16 */
struct _NSZone;
static id 
meth_imp_23(id self, SEL sel, id arg_2, struct _NSZone  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSZone=}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_23(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct _NSZone  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSZone=}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8@12i16 */
static id 
meth_imp_24(id self, SEL sel, id arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_24(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8@12r^f16 */
static id 
meth_imp_25(id self, SEL sel, id arg_2, float  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_25(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	float  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8@12r^{FSRef=[80C]}16 */
struct FSRef {
	unsigned char field_0[80];
};

static id 
meth_imp_26(id self, SEL sel, id arg_2, struct FSRef  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_26(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct FSRef  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8@12r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
struct _NSPoint {
	float field_0;
	float field_1;
};
struct _NSSize {
	float field_0;
	float field_1;
};
struct _NSRect {
	struct _NSPoint field_0;
	struct _NSSize field_1;
};

static id 
meth_imp_27(id self, SEL sel, id arg_2, struct _NSRect  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_27(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct _NSRect  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8@16 */
static id 
meth_imp_28(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_28(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8I12:16 */
static id 
meth_imp_29(id self, SEL sel, unsigned int arg_2, SEL arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_29(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	SEL objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8I12@16 */
static id 
meth_imp_30(id self, SEL sel, unsigned int arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_30(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8I12I16 */
static id 
meth_imp_31(id self, SEL sel, unsigned int arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_31(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8I12^I16 */
static id 
meth_imp_32(id self, SEL sel, unsigned int arg_2, unsigned int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_32(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	unsigned int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8I12^{_NSRange=II}16 */
struct _NSRange {
	unsigned int field_0;
	unsigned int field_1;
};

static id 
meth_imp_33(id self, SEL sel, unsigned int arg_2, struct _NSRange  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_33(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	struct _NSRange  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8L12L16 */
static id 
meth_imp_34(id self, SEL sel, unsigned long arg_2, unsigned long arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("L", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("L", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_34(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned long objc_arg2;
	unsigned long objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("L", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("L", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8Q12 */
static id 
meth_imp_35(id self, SEL sel, unsigned long long arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("Q", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_35(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned long long objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("Q", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8S12@16 */
static id 
meth_imp_36(id self, SEL sel, unsigned short arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_36(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned short objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8S12i16 */
static id 
meth_imp_37(id self, SEL sel, unsigned short arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_37(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned short objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8^?12^v16 */
static id 
meth_imp_38(id self, SEL sel, void*  *arg_2, void  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^?", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_38(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void*  *objc_arg2;
	void  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^?", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8^?12i16 */
static id 
meth_imp_39(id self, SEL sel, void*  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^?", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_39(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void*  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^?", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8^@12@16 */
static id 
meth_imp_40(id self, SEL sel, id  *arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_40(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id  *objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8^@12I16 */
static id 
meth_imp_41(id self, SEL sel, id  *arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_41(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id  *objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8^S12I16 */
static id 
meth_imp_42(id self, SEL sel, unsigned short  *arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_42(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned short  *objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8^i12^i16 */
static id 
meth_imp_43(id self, SEL sel, int  *arg_2, int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_43(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int  *objc_arg2;
	int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8^v12I16 */
static id 
meth_imp_44(id self, SEL sel, void  *arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_44(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void  *objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8^{FSRef=[80C]}12i16 */
static id 
meth_imp_45(id self, SEL sel, struct FSRef  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_45(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct FSRef  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8^{_ProtocolTemplate=#*^{objc_protocol_list}^{objc_method_description_list}^{objc_method_description_list}}12i16 */
struct objc_protocol_list;struct objc_method_description_list;struct objc_method_description_list;struct _ProtocolTemplate {
	Class field_0;
	char* field_1;
	struct objc_protocol_list  *field_2;
	struct objc_method_description_list  *field_3;
	struct objc_method_description_list  *field_4;
};

static id 
meth_imp_46(id self, SEL sel, struct _ProtocolTemplate  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_ProtocolTemplate=#*^{objc_protocol_list=}^{objc_method_description_list=}^{objc_method_description_list=}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_46(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _ProtocolTemplate  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_ProtocolTemplate=#*^{objc_protocol_list=}^{objc_method_description_list=}^{objc_method_description_list=}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8^{hostent=*^*ii^*}12@16 */
struct hostent {
	char* field_0;
	char*  *field_1;
	int field_2;
	int field_3;
	char*  *field_4;
};

static id 
meth_imp_47(id self, SEL sel, struct hostent  *arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{hostent=*^*ii^*}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_47(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct hostent  *objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{hostent=*^*ii^*}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8c12@16 */
static id 
meth_imp_48(id self, SEL sel, char arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_48(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8c12i16 */
static id 
meth_imp_49(id self, SEL sel, char arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_49(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8i12@16 */
static id 
meth_imp_50(id self, SEL sel, int arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_50(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8i12i16 */
static id 
meth_imp_51(id self, SEL sel, int arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_51(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8i12r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
static id 
meth_imp_52(id self, SEL sel, int arg_2, struct _NSRect  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_52(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	struct _NSRect  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8q12 */
static id 
meth_imp_53(id self, SEL sel, long long arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("q", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_53(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	long long objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("q", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8r*12I16 */
static id 
meth_imp_54(id self, SEL sel, char* arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_54(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8r*16 */
static id 
meth_imp_55(id self, SEL sel, char* arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_55(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8r^S12I16 */
static id 
meth_imp_56(id self, SEL sel, unsigned short  *arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_56(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned short  *objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8r^v12I16 */
static id 
meth_imp_57(id self, SEL sel, void  *arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_57(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void  *objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8r^v12r*16 */
static id 
meth_imp_58(id self, SEL sel, void  *arg_2, char* arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_58(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void  *objc_arg2;
	char* objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8r^{_NSSize=ff}12@16 */
static id 
meth_imp_59(id self, SEL sel, struct _NSSize  *arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_59(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSSize  *objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8s12@16 */
static id 
meth_imp_60(id self, SEL sel, short arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_60(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	short objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8{CGPoint=ff}12 */
static id 
meth_imp_61(id self, SEL sel, struct CGPoint arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{CGPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_61(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct CGPoint objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{CGPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8{NSButtonState=iccc}12 */
struct NSButtonState {
	int field_0;
	char field_1;
	char field_2;
	char field_3;
};

static id 
meth_imp_62(id self, SEL sel, struct NSButtonState arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{NSButtonState=iccc}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_62(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct NSButtonState objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{NSButtonState=iccc}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8{_NSPoint=ff}12 */
static id 
meth_imp_63(id self, SEL sel, struct _NSPoint arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_63(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSPoint objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8{_NSRange=II}12 */
static id 
meth_imp_64(id self, SEL sel, struct _NSRange arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_64(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRange objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @12@4:8{_NSSize=ff}12 */
static id 
meth_imp_65(id self, SEL sel, struct _NSSize arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_65(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSSize objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8*12I16c20 */
static id 
meth_imp_66(id self, SEL sel, char* arg_2, unsigned int arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_66(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	unsigned int objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8@12@16c20 */
static id 
meth_imp_67(id self, SEL sel, id arg_2, id arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_67(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8@12^I16c20 */
static id 
meth_imp_68(id self, SEL sel, id arg_2, unsigned int  *arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_68(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	unsigned int  *objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8@12^{?=^SI^SI^SI}16c20 */
static id 
meth_imp_69(id self, SEL sel, id arg_2, struct pyobjcanonymous0  *arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_69(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct pyobjcanonymous0  *objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8@12c16c20 */
static id 
meth_imp_70(id self, SEL sel, id arg_2, char arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_70(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	char objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8^@12c16c20 */
static id 
meth_imp_71(id self, SEL sel, id  *arg_2, char arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_71(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id  *objc_arg2;
	char objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8^S12I16c20 */
static id 
meth_imp_72(id self, SEL sel, unsigned short  *arg_2, unsigned int arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_72(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned short  *objc_arg2;
	unsigned int objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8^{FSRef=[80C]}12c16c20 */
static id 
meth_imp_73(id self, SEL sel, struct FSRef  *arg_2, char arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_73(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct FSRef  *objc_arg2;
	char objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8i12i16c20 */
static id 
meth_imp_74(id self, SEL sel, int arg_2, int arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_74(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	int objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8r^v12I16c20 */
static id 
meth_imp_75(id self, SEL sel, void  *arg_2, unsigned int arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_75(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void  *objc_arg2;
	unsigned int objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8{_NSPoint=ff}12c20 */
static id 
meth_imp_76(id self, SEL sel, struct _NSPoint arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_76(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSPoint objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @13@4:8{_NSRange=II}12c20 */
static id 
meth_imp_77(id self, SEL sel, struct _NSRange arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_77(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRange objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @14@4:8@12@16S20 */
static id 
meth_imp_78(id self, SEL sel, id arg_2, id arg_3, unsigned short arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_78(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	unsigned short objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @14@4:8@12^{tiff=*^{_NXStream}sccsll{?=IIIIIISSSSSSSSSSIIIffSSffII[2S]ISSSSI^S^S^S^S[3^S]*********[2I]II^I^I[2S]^f[2S]S^f^f^f[4^S]S[2S]**I^v}{?=SSL}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}16s20 */
struct _NXStream;struct tiff {
	char* field_0;
	struct _NXStream  *field_1;
	short field_2;
	char field_3;
	char field_4;
	short field_5;
	long field_6;
	long field_7;
	struct pyobjcanonymous0 field_8;
	struct pyobjcanonymous0 field_9;
	int  *field_10;
	int  *field_11;
	int field_12[10];
	long field_13;
	int field_14;
	int field_15;
	long field_16;
	long field_17;
	int field_18;
	long field_19;
	void*  *field_20;
	void*  *field_21;
	void*  *field_22;
	void*  *field_23;
	void*  *field_24;
	void*  *field_25;
	void*  *field_26;
	void*  *field_27;
	void*  *field_28;
	void*  *field_29;
	void*  *field_30;
	void*  *field_31;
	char* field_32;
	int field_33;
	int field_34;
	char* field_35;
	long field_36;
	char* field_37;
	long field_38;
	long field_39;
	int field_40;
	int field_41;
};

static id 
meth_imp_79(id self, SEL sel, id arg_2, struct tiff  *arg_3, short arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{tiff=*^{_NXStream=}sccsll{pyobjcanonymous0=ss}{pyobjcanonymous0=ss}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_79(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct tiff  *objc_arg3;
	short objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{tiff=*^{_NXStream=}sccsll{pyobjcanonymous0=ss}{pyobjcanonymous0=ss}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8*12*20 */
static id 
meth_imp_80(id self, SEL sel, char* arg_2, char* arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_80(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	char* objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8:12@16@20 */
static id 
meth_imp_81(id self, SEL sel, SEL arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_81(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	SEL objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12:16@20 */
static id 
meth_imp_82(id self, SEL sel, id arg_2, SEL arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_82(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	SEL objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12@16*20 */
static id 
meth_imp_83(id self, SEL sel, id arg_2, id arg_3, char* arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_83(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	char* objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12@16@20 */
static id 
meth_imp_84(id self, SEL sel, id arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_84(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12@16I20 */
static id 
meth_imp_85(id self, SEL sel, id arg_2, id arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_85(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12@16^c20 */
static id 
meth_imp_86(id self, SEL sel, id arg_2, id arg_3, char  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_86(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	char  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12@16^{_NSPoint=ff}20 */
static id 
meth_imp_87(id self, SEL sel, id arg_2, id arg_3, struct _NSPoint  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_87(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct _NSPoint  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12@16^{_NSZone=}20 */
struct _NSZone;
static id 
meth_imp_88(id self, SEL sel, id arg_2, id arg_3, struct _NSZone  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSZone=}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_88(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct _NSZone  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSZone=}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12@16i20 */
static id 
meth_imp_89(id self, SEL sel, id arg_2, id arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_89(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12@20 */
static id 
meth_imp_90(id self, SEL sel, id arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_90(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12I16@20 */
static id 
meth_imp_91(id self, SEL sel, id arg_2, unsigned int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_91(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12I16I20 */
static id 
meth_imp_92(id self, SEL sel, id arg_2, unsigned int arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_92(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12I16^{_NSRange=II}20 */
static id 
meth_imp_93(id self, SEL sel, id arg_2, unsigned int arg_3, struct _NSRange  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_93(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	struct _NSRange  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12I16i20 */
static id 
meth_imp_94(id self, SEL sel, id arg_2, unsigned int arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_94(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12^@16^{_NSZone=}20 */
struct _NSZone;
static id 
meth_imp_95(id self, SEL sel, id arg_2, id  *arg_3, struct _NSZone  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSZone=}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_95(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id  *objc_arg3;
	struct _NSZone  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSZone=}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12^{OpaquePMPageFormat=}16^{OpaquePMPrintSettings=}20 */
struct OpaquePMPageFormat;
struct OpaquePMPrintSettings;
static id 
meth_imp_96(id self, SEL sel, id arg_2, struct OpaquePMPageFormat  *arg_3, struct OpaquePMPrintSettings  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{OpaquePMPageFormat=}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{OpaquePMPrintSettings=}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_96(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct OpaquePMPageFormat  *objc_arg3;
	struct OpaquePMPrintSettings  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{OpaquePMPageFormat=}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{OpaquePMPrintSettings=}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12i16:20 */
static id 
meth_imp_97(id self, SEL sel, id arg_2, int arg_3, SEL arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_97(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	int objc_arg3;
	SEL objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12i16@20 */
static id 
meth_imp_98(id self, SEL sel, id arg_2, int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_98(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12i16I20 */
static id 
meth_imp_99(id self, SEL sel, id arg_2, int arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_99(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	int objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12i16i20 */
static id 
meth_imp_100(id self, SEL sel, id arg_2, int arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_100(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	int objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12i16r*20 */
static id 
meth_imp_101(id self, SEL sel, id arg_2, int arg_3, char* arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_101(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	int objc_arg3;
	char* objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12r*16I20 */
static id 
meth_imp_102(id self, SEL sel, id arg_2, char* arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_102(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	char* objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12{_NSPoint=ff}16 */
static id 
meth_imp_103(id self, SEL sel, id arg_2, struct _NSPoint arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_103(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct _NSPoint objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8@12{_NSRange=II}16 */
static id 
meth_imp_104(id self, SEL sel, id arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_104(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8I12^{_NSRange=II}16^I20 */
static id 
meth_imp_105(id self, SEL sel, unsigned int arg_2, struct _NSRange  *arg_3, unsigned int  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_105(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	struct _NSRange  *objc_arg3;
	unsigned int  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8I12r^v16L20 */
static id 
meth_imp_106(id self, SEL sel, unsigned int arg_2, void  *arg_3, unsigned long arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("L", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_106(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	void  *objc_arg3;
	unsigned long objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("L", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8I12{_NSRange=II}16 */
static id 
meth_imp_107(id self, SEL sel, unsigned int arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_107(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8S12I16@20 */
static id 
meth_imp_108(id self, SEL sel, unsigned short arg_2, unsigned int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_108(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned short objc_arg2;
	unsigned int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8S12S16@20 */
static id 
meth_imp_109(id self, SEL sel, unsigned short arg_2, unsigned short arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_109(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned short objc_arg2;
	unsigned short objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8^?12^?16:20 */
static id 
meth_imp_110(id self, SEL sel, void*  *arg_2, void*  *arg_3, SEL arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^?", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^?", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_110(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void*  *objc_arg2;
	void*  *objc_arg3;
	SEL objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^?", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^?", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8^?12^?16I20 */
static id 
meth_imp_111(id self, SEL sel, void*  *arg_2, void*  *arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^?", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^?", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_111(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void*  *objc_arg2;
	void*  *objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^?", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^?", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8^?12^v16@20 */
static id 
meth_imp_112(id self, SEL sel, void*  *arg_2, void  *arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^?", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_112(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void*  *objc_arg2;
	void  *objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^?", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8^@12^@16I20 */
static id 
meth_imp_113(id self, SEL sel, id  *arg_2, id  *arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_113(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id  *objc_arg2;
	id  *objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8^@12^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}20 */
struct _RepresentationInfo;
static id 
meth_imp_114(id self, SEL sel, id  *arg_2, struct _NSRect  *arg_3, struct _RepresentationInfo  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_RepresentationInfo=}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_114(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id  *objc_arg2;
	struct _NSRect  *objc_arg3;
	struct _RepresentationInfo  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_RepresentationInfo=}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12r*16*20 */
static id 
meth_imp_115(id self, SEL sel, struct pyobjcanonymous0  *arg_2, char* arg_3, char* arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_115(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct pyobjcanonymous0  *objc_arg2;
	char* objc_arg3;
	char* objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12r*16r*20 */
static id 
meth_imp_116(id self, SEL sel, struct pyobjcanonymous0  *arg_2, char* arg_3, char* arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_116(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct pyobjcanonymous0  *objc_arg2;
	char* objc_arg3;
	char* objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8i12@16^i20 */
static id 
meth_imp_117(id self, SEL sel, int arg_2, id arg_3, int  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_117(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	id objc_arg3;
	int  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8i12@16i20 */
static id 
meth_imp_118(id self, SEL sel, int arg_2, id arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_118(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	id objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8i12i16@20 */
static id 
meth_imp_119(id self, SEL sel, int arg_2, int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_119(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8i12i16i20 */
static id 
meth_imp_120(id self, SEL sel, int arg_2, int arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_120(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	int objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8i12r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16I20 */
static id 
meth_imp_121(id self, SEL sel, int arg_2, struct _NSRect  *arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_121(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	struct _NSRect  *objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8i12{_NSRange=II}16 */
static id 
meth_imp_122(id self, SEL sel, int arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_122(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8r*12I16I20 */
static id 
meth_imp_123(id self, SEL sel, char* arg_2, unsigned int arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_123(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	unsigned int objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8{_NSRange=II}12^{_NSZone=}20 */
struct _NSZone;
static id 
meth_imp_124(id self, SEL sel, struct _NSRange arg_2, struct _NSZone  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSZone=}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_124(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRange objc_arg2;
	struct _NSZone  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSZone=}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8{_NSSize=ff}12@20 */
static id 
meth_imp_125(id self, SEL sel, struct _NSSize arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_125(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSSize objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @16@4:8{_NSSize=ff}12i20 */
static id 
meth_imp_126(id self, SEL sel, struct _NSSize arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_126(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSSize objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @17@4:8@12@16@20c24 */
static id 
meth_imp_127(id self, SEL sel, id arg_2, id arg_3, id arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_127(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @17@4:8@12@16i20c24 */
static id 
meth_imp_128(id self, SEL sel, id arg_2, id arg_3, int arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_128(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @17@4:8@12^I16I20c24 */
static id 
meth_imp_129(id self, SEL sel, id arg_2, unsigned int  *arg_3, unsigned int arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_129(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	unsigned int  *objc_arg3;
	unsigned int objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @17@4:8I12@16@20c24 */
static id 
meth_imp_130(id self, SEL sel, unsigned int arg_2, id arg_3, id arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_130(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	id objc_arg3;
	id objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @17@4:8Q12s20c24 */
static id 
meth_imp_131(id self, SEL sel, unsigned long long arg_2, short arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("Q", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_131(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned long long objc_arg2;
	short objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("Q", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @17@4:8^{FSCatalogInfo=SsIICCCC{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}[4I][16C][16C]QQQQII}12@16^{FSRef=[80C]}20c24 */
struct UTCDateTime {
	unsigned short field_0;
	unsigned int field_1;
	unsigned short field_2;
};
struct FSCatalogInfo {
	unsigned short field_0;
	short field_1;
	unsigned int field_2;
	unsigned int field_3;
	unsigned char field_4;
	unsigned char field_5;
	unsigned char field_6;
	unsigned char field_7;
	struct UTCDateTime field_8;
	struct UTCDateTime field_9;
	struct UTCDateTime field_10;
	struct UTCDateTime field_11;
	struct UTCDateTime field_12;
	unsigned int field_13[4];
	unsigned char field_14[16];
	unsigned char field_15[16];
	unsigned long long field_16;
	unsigned long long field_17;
	unsigned long long field_18;
	unsigned long long field_19;
	unsigned int field_20;
	unsigned int field_21;
};

static id 
meth_imp_132(id self, SEL sel, struct FSCatalogInfo  *arg_2, id arg_3, struct FSRef  *arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{FSCatalogInfo=SsIICCCC{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}[4I][16C][16C]QQQQII}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_132(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct FSCatalogInfo  *objc_arg2;
	id objc_arg3;
	struct FSRef  *objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{FSCatalogInfo=SsIICCCC{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}[4I][16C][16C]QQQQII}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @17@4:8^{_SelectionAnchor=iii}12^{_SelectionAnchor=iii}16c20c24 */
struct _SelectionAnchor {
	int field_0;
	int field_1;
	int field_2;
};

static id 
meth_imp_133(id self, SEL sel, struct _SelectionAnchor  *arg_2, struct _SelectionAnchor  *arg_3, char arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_SelectionAnchor=iii}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_SelectionAnchor=iii}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_133(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _SelectionAnchor  *objc_arg2;
	struct _SelectionAnchor  *objc_arg3;
	char objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_SelectionAnchor=iii}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_SelectionAnchor=iii}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @17@4:8c12i16i20c24 */
static id 
meth_imp_134(id self, SEL sel, char arg_2, int arg_3, int arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_134(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char objc_arg2;
	int objc_arg3;
	int objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8#12@16@20:24 */
static id 
meth_imp_135(id self, SEL sel, Class arg_2, id arg_3, id arg_4, SEL arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_135(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	Class objc_arg2;
	id objc_arg3;
	id objc_arg4;
	SEL objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8:12i16@20@24 */
static id 
meth_imp_136(id self, SEL sel, SEL arg_2, int arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_136(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	SEL objc_arg2;
	int objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8@12:16@20i24 */
static id 
meth_imp_137(id self, SEL sel, id arg_2, SEL arg_3, id arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_137(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	SEL objc_arg3;
	id objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8@12@16:20@24 */
static id 
meth_imp_138(id self, SEL sel, id arg_2, id arg_3, SEL arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_138(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	SEL objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8@12@16@20@24 */
static id 
meth_imp_139(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_139(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8@12@16@20^@24 */
static id 
meth_imp_140(id self, SEL sel, id arg_2, id arg_3, id arg_4, id  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_140(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8@12@16@20^{_NSZone=}24 */
struct _NSZone;
static id 
meth_imp_141(id self, SEL sel, id arg_2, id arg_3, id arg_4, struct _NSZone  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSZone=}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_141(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct _NSZone  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSZone=}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8@12@16@20i24 */
static id 
meth_imp_142(id self, SEL sel, id arg_2, id arg_3, id arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_142(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8@12@16I20@24 */
static id 
meth_imp_143(id self, SEL sel, id arg_2, id arg_3, unsigned int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_143(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8@12@16c20@24 */
static id 
meth_imp_144(id self, SEL sel, id arg_2, id arg_3, char arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_144(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	char objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8@12@16i20i24 */
static id 
meth_imp_145(id self, SEL sel, id arg_2, id arg_3, int arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_145(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8@12i16i20@24 */
static id 
meth_imp_146(id self, SEL sel, id arg_2, int arg_3, int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_146(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	int objc_arg3;
	int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8@12{_NSRange=II}16i24 */
static id 
meth_imp_147(id self, SEL sel, id arg_2, struct _NSRange arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_147(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct _NSRange objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8I12@16@20^{_NSZone=}24 */
struct _NSZone;
static id 
meth_imp_148(id self, SEL sel, unsigned int arg_2, id arg_3, id arg_4, struct _NSZone  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSZone=}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_148(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct _NSZone  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSZone=}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8I12^{_NSRange=II}16{_NSRange=II}20 */
static id 
meth_imp_149(id self, SEL sel, unsigned int arg_2, struct _NSRange  *arg_3, struct _NSRange arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_149(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	struct _NSRange  *objc_arg3;
	struct _NSRange objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12r*16^*20i24 */
static id 
meth_imp_150(id self, SEL sel, struct pyobjcanonymous0  *arg_2, char* arg_3, char*  *arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^*", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_150(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct pyobjcanonymous0  *objc_arg2;
	char* objc_arg3;
	char*  *objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^*", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8^{__CFSocket=}12i16i20i24 */
struct __CFSocket;
static id 
meth_imp_151(id self, SEL sel, struct __CFSocket  *arg_2, int arg_3, int arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{__CFSocket=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_151(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct __CFSocket  *objc_arg2;
	int objc_arg3;
	int objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{__CFSocket=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8i12i16i20@24 */
static id 
meth_imp_152(id self, SEL sel, int arg_2, int arg_3, int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_152(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	int objc_arg3;
	int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8i12i16i20i24 */
static id 
meth_imp_153(id self, SEL sel, int arg_2, int arg_3, int arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_153(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	int objc_arg3;
	int objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8r*12r*16r*20^{?=b4b1b24(?=*^{?}^{__CFDictionary})}24 */
static id 
meth_imp_154(id self, SEL sel, char* arg_2, char* arg_3, char* arg_4, struct pyobjcanonymous0  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_154(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	char* objc_arg3;
	char* objc_arg4;
	struct pyobjcanonymous0  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8{_NSRange=II}12@20@24 */
static id 
meth_imp_155(id self, SEL sel, struct _NSRange arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_155(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRange objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12 */
static id 
meth_imp_156(id self, SEL sel, struct _NSRect arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_156(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @21@4:8@12@16@20@24c28 */
static id 
meth_imp_157(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_157(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @21@4:8^@12I16@20c24c28 */
static id 
meth_imp_158(id self, SEL sel, id  *arg_2, unsigned int arg_3, id arg_4, char arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_158(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id  *objc_arg2;
	unsigned int objc_arg3;
	id objc_arg4;
	char objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @21@4:8^v12I16c20c24c28 */
static id 
meth_imp_159(id self, SEL sel, void  *arg_2, unsigned int arg_3, char arg_4, char arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_159(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void  *objc_arg2;
	unsigned int objc_arg3;
	char objc_arg4;
	char objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @21@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28 */
static id 
meth_imp_160(id self, SEL sel, struct _NSRect arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_160(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @21@4:8{_NSSize=ff}12i20c24c28 */
static id 
meth_imp_161(id self, SEL sel, struct _NSSize arg_2, int arg_3, char arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_161(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSSize objc_arg2;
	int objc_arg3;
	char objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @22@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12s28 */
static id 
meth_imp_162(id self, SEL sel, struct _NSRect arg_2, short arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_162(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	short objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8*12*16*20*24*28 */
static id 
meth_imp_163(id self, SEL sel, char* arg_2, char* arg_3, char* arg_4, char* arg_5, char* arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_163(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	char* objc_arg3;
	char* objc_arg4;
	char* objc_arg5;
	char* objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8@12@16@20@24@28 */
static id 
meth_imp_164(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_164(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8@12@16@20i24@28 */
static id 
meth_imp_165(id self, SEL sel, id arg_2, id arg_3, id arg_4, int arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_165(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	int objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8@12@16@20{_NSPoint=ff}24 */
static id 
meth_imp_166(id self, SEL sel, id arg_2, id arg_3, id arg_4, struct _NSPoint arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_166(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct _NSPoint objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8@12@16I20@24@28 */
static id 
meth_imp_167(id self, SEL sel, id arg_2, id arg_3, unsigned int arg_4, id arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_167(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	id objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8@12@16{_NSRange=II}20@28 */
static id 
meth_imp_168(id self, SEL sel, id arg_2, id arg_3, struct _NSRange arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_168(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct _NSRange objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8@12I16^{_NSRange=II}20{_NSRange=II}24 */
static id 
meth_imp_169(id self, SEL sel, id arg_2, unsigned int arg_3, struct _NSRange  *arg_4, struct _NSRange arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_169(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	struct _NSRange  *objc_arg4;
	struct _NSRange objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8@12i16{_NSPoint=ff}20^v28 */
static id 
meth_imp_170(id self, SEL sel, id arg_2, int arg_3, struct _NSPoint arg_4, void  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_170(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	int objc_arg3;
	struct _NSPoint objc_arg4;
	void  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
static id 
meth_imp_171(id self, SEL sel, id arg_2, struct _NSRect arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_171(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct _NSRect objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8I12I16@20s24i28 */
static id 
meth_imp_172(id self, SEL sel, unsigned int arg_2, unsigned int arg_3, id arg_4, short arg_5, int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_172(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	unsigned int objc_arg3;
	id objc_arg4;
	short objc_arg5;
	int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8^v12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
static id 
meth_imp_173(id self, SEL sel, void  *arg_2, struct _NSRect arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_173(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void  *objc_arg2;
	struct _NSRect objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8i12@16@20@24i28 */
static id 
meth_imp_174(id self, SEL sel, int arg_2, id arg_3, id arg_4, id arg_5, int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_174(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8i12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
static id 
meth_imp_175(id self, SEL sel, int arg_2, struct _NSRect arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_175(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	struct _NSRect objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I16i20c24@28 */
static id 
meth_imp_176(id self, SEL sel, struct _NSRect  *arg_2, unsigned int arg_3, int arg_4, char arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_176(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect  *objc_arg2;
	unsigned int objc_arg3;
	int objc_arg4;
	char objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8{?=b8b4b1b1b18[8S]}12 */
static id 
meth_imp_177(id self, SEL sel, struct pyobjcanonymous0 arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{pyobjcanonymous0=ss}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_177(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct pyobjcanonymous0 objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{pyobjcanonymous0=ss}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28 */
static id 
meth_imp_178(id self, SEL sel, struct _NSRect arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_178(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @24@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12i28 */
static id 
meth_imp_179(id self, SEL sel, struct _NSRect arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_179(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @25@4:8*12*16*20*24*28c32 */
static id 
meth_imp_180(id self, SEL sel, char* arg_2, char* arg_3, char* arg_4, char* arg_5, char* arg_6, char arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_180(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	char* objc_arg3;
	char* objc_arg4;
	char* objc_arg5;
	char* objc_arg6;
	char objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @25@4:8@12@16@20@24^@28c32 */
static id 
meth_imp_181(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, id  *arg_6, char arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_181(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id  *objc_arg6;
	char objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @25@4:8@12@16i20i24^{_SelectionAnchor=iii}28c32 */
static id 
meth_imp_182(id self, SEL sel, id arg_2, id arg_3, int arg_4, int arg_5, struct _SelectionAnchor  *arg_6, char arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^{_SelectionAnchor=iii}", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_182(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	int objc_arg5;
	struct _SelectionAnchor  *objc_arg6;
	char objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^{_SelectionAnchor=iii}", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @25@4:8i12s16c20c24c28c32 */
static id 
meth_imp_183(id self, SEL sel, int arg_2, short arg_3, char arg_4, char arg_5, char arg_6, char arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_183(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	short objc_arg3;
	char objc_arg4;
	char objc_arg5;
	char objc_arg6;
	char objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @25@4:8{_NSSize=ff}12i20c24c28c32 */
static id 
meth_imp_184(id self, SEL sel, struct _NSSize arg_2, int arg_3, char arg_4, char arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_184(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSSize objc_arg2;
	int objc_arg3;
	char objc_arg4;
	char objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @28@4:8@12@16@20@24@28@32 */
static id 
meth_imp_185(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, id arg_6, id arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_185(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	id objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @28@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32 */
static id 
meth_imp_186(id self, SEL sel, id arg_2, struct _NSRect arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_186(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @28@4:8i12i16i20i24i28i32 */
static id 
meth_imp_187(id self, SEL sel, int arg_2, int arg_3, int arg_4, int arg_5, int arg_6, int arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_187(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	int objc_arg3;
	int objc_arg4;
	int objc_arg5;
	int objc_arg6;
	int objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @28@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I16i20c24@28@32 */
static id 
meth_imp_188(id self, SEL sel, struct _NSRect  *arg_2, unsigned int arg_3, int arg_4, char arg_5, id arg_6, id arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_188(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect  *objc_arg2;
	unsigned int objc_arg3;
	int objc_arg4;
	char objc_arg5;
	id objc_arg6;
	id objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @28@4:8{_NSRange=II}12@20@24{_NSRange=II}28 */
static id 
meth_imp_189(id self, SEL sel, struct _NSRange arg_2, id arg_3, id arg_4, struct _NSRange arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_189(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRange objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct _NSRange objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32 */
static id 
meth_imp_190(id self, SEL sel, struct _NSRect arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_190(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28i32 */
static id 
meth_imp_191(id self, SEL sel, struct _NSRect arg_2, id arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_191(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	id objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I28@32 */
static id 
meth_imp_192(id self, SEL sel, struct _NSRect arg_2, unsigned int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_192(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	unsigned int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8@12@16f36 */
static id 
meth_imp_193(id self, SEL sel, id arg_2, id arg_3, float arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_193(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	float objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8@12I16i20f36 */
static id 
meth_imp_194(id self, SEL sel, id arg_2, unsigned int arg_3, int arg_4, float arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_194(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	int objc_arg4;
	float objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8@12f36 */
static id 
meth_imp_195(id self, SEL sel, id arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_195(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8@12f36@20{_NSPoint=ff}24 */
static id 
meth_imp_196(id self, SEL sel, id arg_2, float arg_3, id arg_4, struct _NSPoint arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_196(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	float objc_arg3;
	id objc_arg4;
	struct _NSPoint objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8@12f36r^f20 */
static id 
meth_imp_197(id self, SEL sel, id arg_2, float arg_3, float  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_197(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	float objc_arg3;
	float  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8@12f36r^f20I24 */
static id 
meth_imp_198(id self, SEL sel, id arg_2, float arg_3, float  *arg_4, unsigned int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_198(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	float objc_arg3;
	float  *objc_arg4;
	unsigned int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8@12f36r^f20i24 */
static id 
meth_imp_199(id self, SEL sel, id arg_2, float arg_3, float  *arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_199(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	float objc_arg3;
	float  *objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8@12i16f36 */
static id 
meth_imp_200(id self, SEL sel, id arg_2, int arg_3, float arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_200(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	int objc_arg3;
	float objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8^{?=*i}12^*16^*20f36 */
static id 
meth_imp_201(id self, SEL sel, struct pyobjcanonymous0  *arg_2, char*  *arg_3, char*  *arg_4, float arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^*", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_201(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct pyobjcanonymous0  *objc_arg2;
	char*  *objc_arg3;
	char*  *objc_arg4;
	float objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^*", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8f36 */
static id 
meth_imp_202(id self, SEL sel, float arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_202(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	float objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8f36@16 */
static id 
meth_imp_203(id self, SEL sel, float arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_203(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	float objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8i12f36 */
static id 
meth_imp_204(id self, SEL sel, int arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_204(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @32@4:8i12f36r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}20r^{_NSPoint=ff}24 */
static id 
meth_imp_205(id self, SEL sel, int arg_2, float arg_3, struct _NSRect  *arg_4, struct _NSPoint  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_205(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	float objc_arg3;
	struct _NSRect  *objc_arg4;
	struct _NSPoint  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8@12:16@20@24@28@32I40 */
static id 
meth_imp_206(id self, SEL sel, id arg_2, SEL arg_3, id arg_4, id arg_5, id arg_6, id arg_7, unsigned int arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_206(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	SEL objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	id objc_arg7;
	unsigned int objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8@12@16c20@24@28:32I40 */
static id 
meth_imp_207(id self, SEL sel, id arg_2, id arg_3, char arg_4, id arg_5, id arg_6, SEL arg_7, unsigned int arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_207(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	id objc_arg3;
	char objc_arg4;
	id objc_arg5;
	id objc_arg6;
	SEL objc_arg7;
	unsigned int objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32@40 */
static id 
meth_imp_208(id self, SEL sel, id arg_2, struct _NSRect arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_208(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8d36 */
static id 
meth_imp_209(id self, SEL sel, double arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_209(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	double objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8d36@20 */
static id 
meth_imp_210(id self, SEL sel, double arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_210(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	double objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8d36@20:24@28c32 */
static id 
meth_imp_211(id self, SEL sel, double arg_2, id arg_3, SEL arg_4, id arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_211(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	double objc_arg2;
	id objc_arg3;
	SEL objc_arg4;
	id objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8d36@20c24 */
static id 
meth_imp_212(id self, SEL sel, double arg_2, id arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_212(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	double objc_arg2;
	id objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8i12@16@20@24@28@32*40 */
static id 
meth_imp_213(id self, SEL sel, int arg_2, id arg_3, id arg_4, id arg_5, id arg_6, id arg_7, char* arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_213(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	id objc_arg7;
	char* objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8i12I16I20I24I28I32@40 */
static id 
meth_imp_214(id self, SEL sel, int arg_2, unsigned int arg_3, unsigned int arg_4, unsigned int arg_5, unsigned int arg_6, unsigned int arg_7, id arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_214(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	unsigned int objc_arg3;
	unsigned int objc_arg4;
	unsigned int objc_arg5;
	unsigned int objc_arg6;
	unsigned int objc_arg7;
	id objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@16@20@24@28i32i40 */
static id 
meth_imp_215(id self, SEL sel, struct _NSRect  *arg_2, id arg_3, id arg_4, id arg_5, id arg_6, int arg_7, int arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_215(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect  *objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	int objc_arg7;
	int objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28I32@40 */
static id 
meth_imp_216(id self, SEL sel, struct _NSRect arg_2, id arg_3, unsigned int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_216(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I28i32c43 */
static id 
meth_imp_217(id self, SEL sel, struct _NSRect arg_2, unsigned int arg_3, int arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_217(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	unsigned int objc_arg3;
	int objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @40@4:8@12d36@24:28@32c43c47 */
static id 
meth_imp_218(id self, SEL sel, id arg_2, double arg_3, id arg_4, SEL arg_5, id arg_6, char arg_7, char arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_218(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	double objc_arg3;
	id objc_arg4;
	SEL objc_arg5;
	id objc_arg6;
	char objc_arg7;
	char objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @40@4:8@12{_NSSize=ff}16f36f44{_NSPoint=ff}36 */
static id 
meth_imp_219(id self, SEL sel, id arg_2, struct _NSSize arg_3, float arg_4, float arg_5, struct _NSPoint arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_219(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct _NSSize objc_arg3;
	float objc_arg4;
	float objc_arg5;
	struct _NSPoint objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @40@4:8f36f44 */
static id 
meth_imp_220(id self, SEL sel, float arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_220(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	float objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @40@4:8f36f44c20 */
static id 
meth_imp_221(id self, SEL sel, float arg_2, float arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_221(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	float objc_arg2;
	float objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I28i32c43@44 */
static id 
meth_imp_222(id self, SEL sel, struct _NSRect arg_2, unsigned int arg_3, int arg_4, char arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_222(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	unsigned int objc_arg3;
	int objc_arg4;
	char objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12i28#32i40i44 */
static id 
meth_imp_223(id self, SEL sel, struct _NSRect arg_2, int arg_3, Class arg_4, int arg_5, int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_223(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	int objc_arg3;
	Class objc_arg4;
	int objc_arg5;
	int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12i28@32i40i44 */
static id 
meth_imp_224(id self, SEL sel, struct _NSRect arg_2, int arg_3, id arg_4, int arg_5, int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_224(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect objc_arg2;
	int objc_arg3;
	id objc_arg4;
	int objc_arg5;
	int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @48@4:8^*12i16i20i24i28c32c43@44i48i52 */
static id 
meth_imp_225(id self, SEL sel, char*  *arg_2, int arg_3, int arg_4, int arg_5, int arg_6, char arg_7, char arg_8, id arg_9, int arg_10, int arg_11)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(11);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_9);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 8, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_10);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 9, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_11);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 10, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_225(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char*  *objc_arg2;
	int objc_arg3;
	int objc_arg4;
	int objc_arg5;
	int objc_arg6;
	char objc_arg7;
	char objc_arg8;
	id objc_arg9;
	int objc_arg10;
	int objc_arg11;
	struct objc_super super;

	if (PyTuple_Size(args) != 10) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 7);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg9);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 8);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg10);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 9);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg11);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8, objc_arg9, objc_arg10, objc_arg11);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @48@4:8i12{_NSPoint=ff}16I24d36i40@44i48i52f44 */
static id 
meth_imp_226(id self, SEL sel, int arg_2, struct _NSPoint arg_3, unsigned int arg_4, double arg_5, int arg_6, id arg_7, int arg_8, int arg_9, float arg_10)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(10);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_9);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 8, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_10);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 9, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_226(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	struct _NSPoint objc_arg3;
	unsigned int objc_arg4;
	double objc_arg5;
	int objc_arg6;
	id objc_arg7;
	int objc_arg8;
	int objc_arg9;
	float objc_arg10;
	struct objc_super super;

	if (PyTuple_Size(args) != 9) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 7);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg9);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 8);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg10);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8, objc_arg9, objc_arg10);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @4@4:8 */
static id 
meth_imp_227(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_227(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @52@4:8i12{_NSPoint=ff}16I24d36i40@44i48i52^v56 */
static id 
meth_imp_228(id self, SEL sel, int arg_2, struct _NSPoint arg_3, unsigned int arg_4, double arg_5, int arg_6, id arg_7, int arg_8, int arg_9, void  *arg_10)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(10);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_9);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 8, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_10);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 9, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_228(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	struct _NSPoint objc_arg3;
	unsigned int objc_arg4;
	double objc_arg5;
	int objc_arg6;
	id objc_arg7;
	int objc_arg8;
	int objc_arg9;
	void  *objc_arg10;
	struct objc_super super;

	if (PyTuple_Size(args) != 9) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 7);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg9);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 8);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg10);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8, objc_arg9, objc_arg10);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @52@4:8i12{_NSPoint=ff}16I24d36i40@44s50i52i56 */
static id 
meth_imp_229(id self, SEL sel, int arg_2, struct _NSPoint arg_3, unsigned int arg_4, double arg_5, int arg_6, id arg_7, short arg_8, int arg_9, int arg_10)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(10);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_9);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 8, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_10);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 9, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_229(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	struct _NSPoint objc_arg3;
	unsigned int objc_arg4;
	double objc_arg5;
	int objc_arg6;
	id objc_arg7;
	short objc_arg8;
	int objc_arg9;
	int objc_arg10;
	struct objc_super super;

	if (PyTuple_Size(args) != 9) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 7);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg9);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 8);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg10);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8, objc_arg9, objc_arg10);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @56@4:8^*12i16i20i24i28c32c43@44i48i52{_NSSize=ff}56 */
static id 
meth_imp_230(id self, SEL sel, char*  *arg_2, int arg_3, int arg_4, int arg_5, int arg_6, char arg_7, char arg_8, id arg_9, int arg_10, int arg_11, struct _NSSize arg_12)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(12);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_9);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 8, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_10);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 9, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_11);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 10, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_12);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 11, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_230(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char*  *objc_arg2;
	int objc_arg3;
	int objc_arg4;
	int objc_arg5;
	int objc_arg6;
	char objc_arg7;
	char objc_arg8;
	id objc_arg9;
	int objc_arg10;
	int objc_arg11;
	struct _NSSize objc_arg12;
	struct objc_super super;

	if (PyTuple_Size(args) != 11) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 7);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg9);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 8);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg10);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 9);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg11);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 10);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg12);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8, objc_arg9, objc_arg10, objc_arg11, objc_arg12);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @56@4:8f36f44f52f60 */
static id 
meth_imp_231(id self, SEL sel, float arg_2, float arg_3, float arg_4, float arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_231(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	float objc_arg2;
	float objc_arg3;
	float objc_arg4;
	float objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @56@4:8i12{_NSPoint=ff}16I24d36i40@44@48@52c59S62 */
static id 
meth_imp_232(id self, SEL sel, int arg_2, struct _NSPoint arg_3, unsigned int arg_4, double arg_5, int arg_6, id arg_7, id arg_8, id arg_9, char arg_10, unsigned short arg_11)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(11);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_9);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 8, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_10);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 9, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_11);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 10, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_232(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	struct _NSPoint objc_arg3;
	unsigned int objc_arg4;
	double objc_arg5;
	int objc_arg6;
	id objc_arg7;
	id objc_arg8;
	id objc_arg9;
	char objc_arg10;
	unsigned short objc_arg11;
	struct objc_super super;

	if (PyTuple_Size(args) != 10) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 7);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg9);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 8);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg10);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 9);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg11);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8, objc_arg9, objc_arg10, objc_arg11);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @5@4:8C12 */
static id 
meth_imp_233(id self, SEL sel, unsigned char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("C", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_233(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("C", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @5@4:8c12 */
static id 
meth_imp_234(id self, SEL sel, char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_234(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @64@4:8f36f44f52f60f68 */
static id 
meth_imp_235(id self, SEL sel, float arg_2, float arg_3, float arg_4, float arg_5, float arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_235(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	float objc_arg2;
	float objc_arg3;
	float objc_arg4;
	float objc_arg5;
	float objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @6@4:8S12 */
static id 
meth_imp_236(id self, SEL sel, unsigned short arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_236(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned short objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @6@4:8s12 */
static id 
meth_imp_237(id self, SEL sel, short arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_237(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	short objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8#12 */
static id 
meth_imp_238(id self, SEL sel, Class arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_238(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	Class objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8*12 */
static id 
meth_imp_239(id self, SEL sel, char* arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_239(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8:12 */
static id 
meth_imp_240(id self, SEL sel, SEL arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_240(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	SEL objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8@12 */
static id 
meth_imp_241(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_241(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8I12 */
static id 
meth_imp_242(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_242(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8L12 */
static id 
meth_imp_243(id self, SEL sel, unsigned long arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("L", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_243(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned long objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("L", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^c12 */
static id 
meth_imp_244(id self, SEL sel, char  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_244(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^i12 */
static id 
meth_imp_245(id self, SEL sel, int  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_245(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^v12 */
static id 
meth_imp_246(id self, SEL sel, void  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_246(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12 */
static id 
meth_imp_247(id self, SEL sel, struct pyobjcanonymous0  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_247(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct pyobjcanonymous0  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{FSRef=[80C]}12 */
static id 
meth_imp_248(id self, SEL sel, struct FSRef  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_248(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct FSRef  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{NSCharSetPrivateStruct=i[4i]iiii[1i]}12 */
struct NSCharSetPrivateStruct {
	int field_0;
	int field_1[4];
	int field_2;
	int field_3;
	int field_4;
	int field_5;
	int field_6[1];
};

static id 
meth_imp_249(id self, SEL sel, struct NSCharSetPrivateStruct  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{NSCharSetPrivateStruct=i[4i]iiii[1i]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_249(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct NSCharSetPrivateStruct  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{NSCharSetPrivateStruct=i[4i]iiii[1i]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{_NSPoint=ff}12 */
static id 
meth_imp_250(id self, SEL sel, struct _NSPoint  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_250(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSPoint  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12 */
static id 
meth_imp_251(id self, SEL sel, struct _NSRect  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_251(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{_NSRefCountedRunArray=IIIIII[0{_NSRunArrayItem=I@}]}12 */
struct _NSRunArrayItem {
	unsigned int field_0;
	id field_1;
};
struct _NSRefCountedRunArray {
	unsigned int field_0;
	unsigned int field_1;
	unsigned int field_2;
	unsigned int field_3;
	unsigned int field_4;
	unsigned int field_5;
	struct _NSRunArrayItem field_6[0];
};

static id 
meth_imp_252(id self, SEL sel, struct _NSRefCountedRunArray  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRefCountedRunArray=IIIIII[0{_NSRunArrayItem=I@}]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_252(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRefCountedRunArray  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRefCountedRunArray=IIIIII[0{_NSRunArrayItem=I@}]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{_NSRulebookSetHeader=i[4L]iiii[1i]}12 */
struct _NSRulebookSetHeader {
	int field_0;
	unsigned long field_1[4];
	int field_2;
	int field_3;
	int field_4;
	int field_5;
	int field_6[1];
};

static id 
meth_imp_253(id self, SEL sel, struct _NSRulebookSetHeader  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRulebookSetHeader=i[4L]iiii[1i]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_253(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRulebookSetHeader  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRulebookSetHeader=i[4L]iiii[1i]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{_NSSize=ff}12 */
static id 
meth_imp_254(id self, SEL sel, struct _NSSize  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_254(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSSize  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{_NSStringBuffer=II@II[32S]S}12 */
struct _NSStringBuffer {
	unsigned int field_0;
	unsigned int field_1;
	id field_2;
	unsigned int field_3;
	unsigned int field_4;
	unsigned short field_5[32];
	unsigned short field_6;
};

static id 
meth_imp_255(id self, SEL sel, struct _NSStringBuffer  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSStringBuffer=II@II[32S]S}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_255(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSStringBuffer  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSStringBuffer=II@II[32S]S}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{_NSZone=}12 */
struct _NSZone;
static id 
meth_imp_256(id self, SEL sel, struct _NSZone  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSZone=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_256(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSZone  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSZone=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}12 */
struct _RepresentationInfo;
static id 
meth_imp_257(id self, SEL sel, struct _RepresentationInfo  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_RepresentationInfo=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_257(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _RepresentationInfo  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_RepresentationInfo=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{__CFNotificationCenter=}12 */
struct __CFNotificationCenter;
static id 
meth_imp_258(id self, SEL sel, struct __CFNotificationCenter  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{__CFNotificationCenter=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_258(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct __CFNotificationCenter  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{__CFNotificationCenter=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{_object=i^{_typeobject}}12 */
static id 
meth_imp_259(id self, SEL sel, struct _object  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_object=i^{_typeobject=}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_259(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _object  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_object=i^{_typeobject=}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{hostent=*^*ii^*}12 */
static id 
meth_imp_260(id self, SEL sel, struct hostent  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{hostent=*^*ii^*}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_260(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct hostent  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{hostent=*^*ii^*}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8^{stat=iISSIIi{timespec=ii}{timespec=ii}{timespec=ii}qqIIIi[2q]}12 */
static id 
meth_imp_261(id self, SEL sel, struct stat  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{stat=iISSIIi{timespec=ii}{timespec=ii}{timespec=ii}qqIIIi[2q]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_261(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct stat  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{stat=iISSIIi{timespec=ii}{timespec=ii}{timespec=ii}qqIIIi[2q]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8i12 */
static id 
meth_imp_262(id self, SEL sel, int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_262(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8l12 */
static id 
meth_imp_263(id self, SEL sel, long arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("l", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_263(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	long objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("l", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8r*12 */
static id 
meth_imp_264(id self, SEL sel, char* arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_264(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char* objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8r^v12 */
static id 
meth_imp_265(id self, SEL sel, void  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_265(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8r^{FSRef=[80C]}12 */
static id 
meth_imp_266(id self, SEL sel, struct FSRef  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_266(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct FSRef  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @8@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12 */
static id 
meth_imp_267(id self, SEL sel, struct _NSRect  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_267(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _NSRect  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @9@4:8:12c16 */
static id 
meth_imp_268(id self, SEL sel, SEL arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_268(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	SEL objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @9@4:8@12c16 */
static id 
meth_imp_269(id self, SEL sel, id arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_269(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @9@4:8I12c16 */
static id 
meth_imp_270(id self, SEL sel, unsigned int arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_270(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	unsigned int objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @9@4:8^@12c16 */
static id 
meth_imp_271(id self, SEL sel, id  *arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_271(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	id  *objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @9@4:8^v12c16 */
static id 
meth_imp_272(id self, SEL sel, void  *arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_272(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	void  *objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @9@4:8^{OpaqueWindowPtr=}12c16 */
struct OpaqueWindowPtr;
static id 
meth_imp_273(id self, SEL sel, struct OpaqueWindowPtr  *arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{OpaqueWindowPtr=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_273(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct OpaqueWindowPtr  *objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{OpaqueWindowPtr=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @9@4:8^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}12c16 */
struct _RepresentationInfo;
static id 
meth_imp_274(id self, SEL sel, struct _RepresentationInfo  *arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_RepresentationInfo=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_274(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _RepresentationInfo  *objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_RepresentationInfo=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @9@4:8^{_SelectionAnchor=iii}12c16 */
static id 
meth_imp_275(id self, SEL sel, struct _SelectionAnchor  *arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_SelectionAnchor=iii}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_275(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	struct _SelectionAnchor  *objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_SelectionAnchor=iii}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @9@4:8c12c16 */
static id 
meth_imp_276(id self, SEL sel, char arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_276(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	char objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: @9@4:8i12c16 */
static id 
meth_imp_277(id self, SEL sel, int arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	id objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("@", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_277(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_retval;
	int objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (id)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("@", &objc_retval);
	return v;
}


/* signature: C14@4:8I12^{OpaqueMenuHandle=}16S20 */
struct OpaqueMenuHandle;
static unsigned char 
meth_imp_278(id self, SEL sel, unsigned int arg_2, struct OpaqueMenuHandle  *arg_3, unsigned short arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{OpaqueMenuHandle=}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("C", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_278(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned char objc_retval;
	unsigned int objc_arg2;
	struct OpaqueMenuHandle  *objc_arg3;
	unsigned short objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{OpaqueMenuHandle=}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("C", &objc_retval);
	return v;
}


/* signature: C4@4:8 */
static unsigned char 
meth_imp_279(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned char objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("C", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_279(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned char objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (unsigned char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("C", &objc_retval);
	return v;
}


/* signature: I12@4:8:12@16 */
static unsigned int 
meth_imp_280(id self, SEL sel, SEL arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_280(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	SEL objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I12@4:8@12@16 */
static unsigned int 
meth_imp_281(id self, SEL sel, id arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_281(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I12@4:8@12I16 */
static unsigned int 
meth_imp_282(id self, SEL sel, id arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_282(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I12@4:8I12*16 */
static unsigned int 
meth_imp_283(id self, SEL sel, unsigned int arg_2, char* arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_283(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	unsigned int objc_arg2;
	char* objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I12@4:8I12^c16 */
static unsigned int 
meth_imp_284(id self, SEL sel, unsigned int arg_2, char  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_284(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	unsigned int objc_arg2;
	char  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I12@4:8^I12@16 */
static unsigned int 
meth_imp_285(id self, SEL sel, unsigned int  *arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_285(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	unsigned int  *objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I12@4:8r^v12I16 */
static unsigned int 
meth_imp_286(id self, SEL sel, void  *arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_286(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	void  *objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I12@4:8{_NSPoint=ff}12 */
static unsigned int 
meth_imp_287(id self, SEL sel, struct _NSPoint arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_287(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	struct _NSPoint objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I13@4:8@12@16c20 */
static unsigned int 
meth_imp_288(id self, SEL sel, id arg_2, id arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_288(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	id objc_arg2;
	id objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I16@4:8@12@16@20 */
static unsigned int 
meth_imp_289(id self, SEL sel, id arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_289(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I16@4:8@12{_NSRange=II}16 */
static unsigned int 
meth_imp_290(id self, SEL sel, id arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_290(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	id objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I16@4:8^I12@16I20 */
static unsigned int 
meth_imp_291(id self, SEL sel, unsigned int  *arg_2, id arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_291(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	unsigned int  *objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I16@4:8^I12{_NSRange=II}16 */
static unsigned int 
meth_imp_292(id self, SEL sel, unsigned int  *arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_292(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	unsigned int  *objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I16@4:8{_NSPoint=ff}12@20 */
static unsigned int 
meth_imp_293(id self, SEL sel, struct _NSPoint arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_293(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	struct _NSPoint objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I17@4:8@12i16@20c24 */
static unsigned int 
meth_imp_294(id self, SEL sel, id arg_2, int arg_3, id arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_294(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	id objc_arg2;
	int objc_arg3;
	id objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I17@4:8@12{_NSRange=II}16c24 */
static unsigned int 
meth_imp_295(id self, SEL sel, id arg_2, struct _NSRange arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_295(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	id objc_arg2;
	struct _NSRange objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I20@4:8^@12c16^@20@24 */
static unsigned int 
meth_imp_296(id self, SEL sel, id  *arg_2, char arg_3, id  *arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_296(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	id  *objc_arg2;
	char objc_arg3;
	id  *objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I20@4:8{_NSPoint=ff}12@20^f24 */
static unsigned int 
meth_imp_297(id self, SEL sel, struct _NSPoint arg_2, id arg_3, float  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_297(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	struct _NSPoint objc_arg2;
	id objc_arg3;
	float  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I24@4:8@12I16{_NSRange=II}20@28 */
static unsigned int 
meth_imp_298(id self, SEL sel, id arg_2, unsigned int arg_3, struct _NSRange arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_298(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	struct _NSRange objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I28@4:8{_NSRange=II}12^I20^I24^i28^c32 */
static unsigned int 
meth_imp_299(id self, SEL sel, struct _NSRange arg_2, unsigned int  *arg_3, unsigned int  *arg_4, int  *arg_5, char  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_299(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	struct _NSRange objc_arg2;
	unsigned int  *objc_arg3;
	unsigned int  *objc_arg4;
	int  *objc_arg5;
	char  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I4@4:8 */
static unsigned int 
meth_imp_300(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_300(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I5@4:8c12 */
static unsigned int 
meth_imp_301(id self, SEL sel, char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_301(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I6@4:8S12 */
static unsigned int 
meth_imp_302(id self, SEL sel, unsigned short arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_302(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	unsigned short objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I8@4:8:12 */
static unsigned int 
meth_imp_303(id self, SEL sel, SEL arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_303(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	SEL objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I8@4:8@12 */
static unsigned int 
meth_imp_304(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_304(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I8@4:8I12 */
static unsigned int 
meth_imp_305(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_305(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I8@4:8^I12 */
static unsigned int 
meth_imp_306(id self, SEL sel, unsigned int  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_306(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	unsigned int  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I8@4:8^i12 */
static unsigned int 
meth_imp_307(id self, SEL sel, int  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_307(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	int  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I8@4:8i12 */
static unsigned int 
meth_imp_308(id self, SEL sel, int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_308(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I8@4:8l12 */
static unsigned int 
meth_imp_309(id self, SEL sel, long arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("l", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_309(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	long objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("l", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: I9@4:8I12c16 */
static unsigned int 
meth_imp_310(id self, SEL sel, unsigned int arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_310(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_retval;
	unsigned int objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("I", &objc_retval);
	return v;
}


/* signature: L4@4:8 */
static unsigned long 
meth_imp_311(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned long objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("L", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_311(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned long objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (unsigned long)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("L", &objc_retval);
	return v;
}


/* signature: L8@4:8@12 */
static unsigned long 
meth_imp_312(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned long objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("L", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_312(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned long objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned long)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("L", &objc_retval);
	return v;
}


/* signature: S4@4:8 */
static unsigned short 
meth_imp_313(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned short objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("S", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_313(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned short objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (unsigned short)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("S", &objc_retval);
	return v;
}


/* signature: S8@4:8I12 */
static unsigned short 
meth_imp_314(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned short objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("S", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_314(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned short objc_retval;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (unsigned short)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("S", &objc_retval);
	return v;
}


/* signature: ^*4@4:8 */
static char*  *
meth_imp_315(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char*  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^*", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_315(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char*  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (char*  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^*", &objc_retval);
	return v;
}


/* signature: ^?8@4:8:12 */
static void*  *
meth_imp_316(id self, SEL sel, SEL arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	void*  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^?", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_316(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void*  *objc_retval;
	SEL objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (void*  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^?", &objc_retval);
	return v;
}


/* signature: ^S4@4:8 */
static unsigned short  *
meth_imp_317(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned short  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^S", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_317(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned short  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (unsigned short  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^S", &objc_retval);
	return v;
}


/* signature: ^i12@4:8@12^i16 */
static int  *
meth_imp_318(id self, SEL sel, id arg_2, int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int  *objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_318(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_retval;
	id objc_arg2;
	int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^i", &objc_retval);
	return v;
}


/* signature: ^i4@4:8 */
static int  *
meth_imp_319(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_319(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (int  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^i", &objc_retval);
	return v;
}


/* signature: ^i6@4:8S12 */
static int  *
meth_imp_320(id self, SEL sel, unsigned short arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_320(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_retval;
	unsigned short objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^i", &objc_retval);
	return v;
}


/* signature: ^v12@4:8I12^{_NSRange=II}16 */
static void  *
meth_imp_321(id self, SEL sel, unsigned int arg_2, struct _NSRange  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	void  *objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^v", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_321(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_retval;
	unsigned int objc_arg2;
	struct _NSRange  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (void  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^v", &objc_retval);
	return v;
}


/* signature: ^v20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12 */
static void  *
meth_imp_322(id self, SEL sel, struct _NSRect arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	void  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^v", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_322(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_retval;
	struct _NSRect objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (void  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^v", &objc_retval);
	return v;
}


/* signature: ^v4@4:8 */
static void  *
meth_imp_323(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	void  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^v", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_323(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (void  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^v", &objc_retval);
	return v;
}


/* signature: ^v5@4:8c12 */
static void  *
meth_imp_324(id self, SEL sel, char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	void  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^v", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_324(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_retval;
	char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (void  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^v", &objc_retval);
	return v;
}


/* signature: ^v8@4:8@12 */
static void  *
meth_imp_325(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	void  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^v", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_325(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (void  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^v", &objc_retval);
	return v;
}


/* signature: ^v8@4:8I12 */
static void  *
meth_imp_326(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	void  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^v", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_326(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_retval;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (void  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^v", &objc_retval);
	return v;
}


/* signature: ^v8@4:8^I12 */
static void  *
meth_imp_327(id self, SEL sel, unsigned int  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	void  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^v", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_327(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_retval;
	unsigned int  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (void  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^v", &objc_retval);
	return v;
}


/* signature: ^{?=^{OpaquePMPrintSession}^{OpaquePMPrintSettings}^{OpaquePMPageFormat}}4@4:8 */
static struct pyobjcanonymous0  *
meth_imp_328(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct pyobjcanonymous0  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_328(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct pyobjcanonymous0  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct pyobjcanonymous0  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &objc_retval);
	return v;
}


/* signature: ^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12@4:8r*12^{?=b4b1b24(?=*^{?}^{__CFDictionary})}16 */
static struct pyobjcanonymous0  *
meth_imp_329(id self, SEL sel, char* arg_2, struct pyobjcanonymous0  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct pyobjcanonymous0  *objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_329(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct pyobjcanonymous0  *objc_retval;
	char* objc_arg2;
	struct pyobjcanonymous0  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct pyobjcanonymous0  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &objc_retval);
	return v;
}


/* signature: ^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12@4:8r*12r*16 */
static struct pyobjcanonymous0  *
meth_imp_330(id self, SEL sel, char* arg_2, char* arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct pyobjcanonymous0  *objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_330(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct pyobjcanonymous0  *objc_retval;
	char* objc_arg2;
	char* objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct pyobjcanonymous0  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &objc_retval);
	return v;
}


/* signature: ^{?=b4b1b24(?=*^{?}^{__CFDictionary})}8@4:8i12 */
static struct pyobjcanonymous0  *
meth_imp_331(id self, SEL sel, int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct pyobjcanonymous0  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_331(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct pyobjcanonymous0  *objc_retval;
	int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct pyobjcanonymous0  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &objc_retval);
	return v;
}


/* signature: ^{AEDesc=I^^{OpaqueAEDataStorageType}}4@4:8 */
struct OpaqueAEDataStorageType;struct AEDesc {
	unsigned int field_0;
	struct OpaqueAEDataStorageType  * *field_1;
};

static struct AEDesc  *
meth_imp_332(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct AEDesc  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{AEDesc=I^^{OpaqueAEDataStorageType=}}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_332(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct AEDesc  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct AEDesc  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{AEDesc=I^^{OpaqueAEDataStorageType=}}", &objc_retval);
	return v;
}


/* signature: ^{CGFont=^{CGFontVTable}Ii^{CGEncoding}^{CGCMap}^{CGAdvanceSet}^{CGAdvanceSet}i^{CGFontCache}^vb1b1b1b1}4@4:8 */
struct CGFontVTable;struct CGEncoding;struct CGCMap;struct CGAdvanceSet;struct CGAdvanceSet;struct CGFontCache;struct CGFont {
	struct CGFontVTable  *field_0;
	unsigned int field_1;
	int field_2;
	struct CGEncoding  *field_3;
	struct CGCMap  *field_4;
	struct CGAdvanceSet  *field_5;
	struct CGAdvanceSet  *field_6;
	int field_7;
	struct CGFontCache  *field_8;
	void  *field_9;
	int field_10:1;
	int field_11:1;
	int field_12:1;
	int field_13:1;
};

static struct CGFont  *
meth_imp_333(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct CGFont  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{CGFont=^{CGFontVTable=}Ii^{CGEncoding=}^{CGCMap=}^{CGAdvanceSet=}^{CGAdvanceSet=}i^{CGFontCache=}^vb1b1b1b1}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_333(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct CGFont  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct CGFont  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{CGFont=^{CGFontVTable=}Ii^{CGEncoding=}^{CGCMap=}^{CGAdvanceSet=}^{CGAdvanceSet=}i^{CGFontCache=}^vb1b1b1b1}", &objc_retval);
	return v;
}


/* signature: ^{CGPDFDocument=}4@4:8 */
struct CGPDFDocument;
static struct CGPDFDocument  *
meth_imp_334(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct CGPDFDocument  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{CGPDFDocument=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_334(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct CGPDFDocument  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct CGPDFDocument  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{CGPDFDocument=}", &objc_retval);
	return v;
}


/* signature: ^{ComponentInstanceRecord=[1l]}5@4:8c12 */
struct ComponentInstanceRecord {
	long field_0[1];
};

static struct ComponentInstanceRecord  *
meth_imp_335(id self, SEL sel, char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct ComponentInstanceRecord  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{ComponentInstanceRecord=[1l]}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_335(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct ComponentInstanceRecord  *objc_retval;
	char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct ComponentInstanceRecord  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{ComponentInstanceRecord=[1l]}", &objc_retval);
	return v;
}


/* signature: ^{FSRef=[80C]}4@4:8 */
static struct FSRef  *
meth_imp_336(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct FSRef  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_336(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct FSRef  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct FSRef  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{FSRef=[80C]}", &objc_retval);
	return v;
}


/* signature: ^{OpaqueCoreDragHandler=}4@4:8 */
struct OpaqueCoreDragHandler;
static struct OpaqueCoreDragHandler  *
meth_imp_337(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct OpaqueCoreDragHandler  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{OpaqueCoreDragHandler=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_337(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaqueCoreDragHandler  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct OpaqueCoreDragHandler  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{OpaqueCoreDragHandler=}", &objc_retval);
	return v;
}


/* signature: ^{OpaqueGrafPtr=}4@4:8 */
struct OpaqueGrafPtr;
static struct OpaqueGrafPtr  *
meth_imp_338(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct OpaqueGrafPtr  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{OpaqueGrafPtr=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_338(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaqueGrafPtr  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct OpaqueGrafPtr  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{OpaqueGrafPtr=}", &objc_retval);
	return v;
}


/* signature: ^{OpaqueIconRef=}4@4:8 */
struct OpaqueIconRef;
static struct OpaqueIconRef  *
meth_imp_339(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct OpaqueIconRef  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{OpaqueIconRef=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_339(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaqueIconRef  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct OpaqueIconRef  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{OpaqueIconRef=}", &objc_retval);
	return v;
}


/* signature: ^{OpaquePMPageFormat=}4@4:8 */
struct OpaquePMPageFormat;
static struct OpaquePMPageFormat  *
meth_imp_340(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct OpaquePMPageFormat  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{OpaquePMPageFormat=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_340(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaquePMPageFormat  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct OpaquePMPageFormat  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{OpaquePMPageFormat=}", &objc_retval);
	return v;
}


/* signature: ^{OpaquePMPrintSession=}4@4:8 */
struct OpaquePMPrintSession;
static struct OpaquePMPrintSession  *
meth_imp_341(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct OpaquePMPrintSession  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{OpaquePMPrintSession=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_341(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaquePMPrintSession  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct OpaquePMPrintSession  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{OpaquePMPrintSession=}", &objc_retval);
	return v;
}


/* signature: ^{OpaquePMPrintSettings=}4@4:8 */
struct OpaquePMPrintSettings;
static struct OpaquePMPrintSettings  *
meth_imp_342(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct OpaquePMPrintSettings  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{OpaquePMPrintSettings=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_342(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaquePMPrintSettings  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct OpaquePMPrintSettings  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{OpaquePMPrintSettings=}", &objc_retval);
	return v;
}


/* signature: ^{OpaqueWindowPtr=}4@4:8 */
struct OpaqueWindowPtr;
static struct OpaqueWindowPtr  *
meth_imp_343(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct OpaqueWindowPtr  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{OpaqueWindowPtr=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_343(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaqueWindowPtr  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct OpaqueWindowPtr  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{OpaqueWindowPtr=}", &objc_retval);
	return v;
}


/* signature: ^{_CoercerData=@:}12@4:8#12#16 */
struct _CoercerData {
	id field_0;
	SEL field_1;
};

static struct _CoercerData  *
meth_imp_344(id self, SEL sel, Class arg_2, Class arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _CoercerData  *objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_CoercerData=@:}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_344(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _CoercerData  *objc_retval;
	Class objc_arg2;
	Class objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _CoercerData  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_CoercerData=@:}", &objc_retval);
	return v;
}


/* signature: ^{_NSFaceInfo=i^{_NSFaceInfo}@i{_NSFont_faceFlags=b1b1b1b1b1b1b1b1b1b1b22}^{_NSFontMetrics}^{_NSCGSFontMetrics}}8@4:8^{_NSFaceInfo=i^{_NSFaceInfo}@i{_NSFont_faceFlags=b1b1b1b1b1b1b1b1b1b1b22}^{_NSFontMetrics}^{_NSCGSFontMetrics}}12 */
struct _NSFaceInfo;
struct _NSFaceInfo;
static struct _NSFaceInfo  *
meth_imp_345(id self, SEL sel, struct _NSFaceInfo  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSFaceInfo  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSFaceInfo=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSFaceInfo=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_345(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSFaceInfo  *objc_retval;
	struct _NSFaceInfo  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSFaceInfo=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _NSFaceInfo  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSFaceInfo=}", &objc_retval);
	return v;
}


/* signature: ^{_NSMapTable=}5@4:8c12 */
struct _NSMapTable;
static struct _NSMapTable  *
meth_imp_346(id self, SEL sel, char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSMapTable  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSMapTable=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_346(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSMapTable  *objc_retval;
	char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _NSMapTable  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSMapTable=}", &objc_retval);
	return v;
}


/* signature: ^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}12@4:8@12@16 */
struct _NSModalSession;
static struct _NSModalSession  *
meth_imp_347(id self, SEL sel, id arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSModalSession  *objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSModalSession=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_347(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSModalSession  *objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _NSModalSession  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSModalSession=}", &objc_retval);
	return v;
}


/* signature: ^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}24@4:8@12@16@20:24^v28 */
struct _NSModalSession;
static struct _NSModalSession  *
meth_imp_348(id self, SEL sel, id arg_2, id arg_3, id arg_4, SEL arg_5, void  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSModalSession  *objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSModalSession=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_348(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSModalSession  *objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	SEL objc_arg5;
	void  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _NSModalSession  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSModalSession=}", &objc_retval);
	return v;
}


/* signature: ^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}8@4:8@12 */
struct _NSModalSession;
static struct _NSModalSession  *
meth_imp_349(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSModalSession  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSModalSession=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_349(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSModalSession  *objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _NSModalSession  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSModalSession=}", &objc_retval);
	return v;
}


/* signature: ^{_NSRect={_NSPoint=ff}{_NSSize=ff}}20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12 */
static struct _NSRect  *
meth_imp_350(id self, SEL sel, struct _NSRect arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSRect  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_350(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect  *objc_retval;
	struct _NSRect objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _NSRect  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &objc_retval);
	return v;
}


/* signature: ^{_NSRect={_NSPoint=ff}{_NSSize=ff}}28@4:8{_NSRange=II}12{_NSRange=II}20@28^I32 */
static struct _NSRect  *
meth_imp_351(id self, SEL sel, struct _NSRange arg_2, struct _NSRange arg_3, id arg_4, unsigned int  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSRect  *objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_351(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect  *objc_retval;
	struct _NSRange objc_arg2;
	struct _NSRange objc_arg3;
	id objc_arg4;
	unsigned int  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _NSRect  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &objc_retval);
	return v;
}


/* signature: ^{_NSRulebookSetHeader=i[4L]iiii[1i]}4@4:8 */
static struct _NSRulebookSetHeader  *
meth_imp_352(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSRulebookSetHeader  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSRulebookSetHeader=i[4L]iiii[1i]}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_352(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRulebookSetHeader  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct _NSRulebookSetHeader  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSRulebookSetHeader=i[4L]iiii[1i]}", &objc_retval);
	return v;
}


/* signature: ^{_NSRulebookSetHeader=i[4L]iiii[1i]}8@4:8I12 */
static struct _NSRulebookSetHeader  *
meth_imp_353(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSRulebookSetHeader  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSRulebookSetHeader=i[4L]iiii[1i]}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_353(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRulebookSetHeader  *objc_retval;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _NSRulebookSetHeader  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSRulebookSetHeader=i[4L]iiii[1i]}", &objc_retval);
	return v;
}


/* signature: ^{_NSRulebookTestStruct=iii[12i]}8@4:8I12 */
struct _NSRulebookTestStruct {
	int field_0;
	int field_1;
	int field_2;
	int field_3[12];
};

static struct _NSRulebookTestStruct  *
meth_imp_354(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSRulebookTestStruct  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSRulebookTestStruct=iii[12i]}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_354(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRulebookTestStruct  *objc_retval;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _NSRulebookTestStruct  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSRulebookTestStruct=iii[12i]}", &objc_retval);
	return v;
}


/* signature: ^{_NSTypesetterGlyphInfo={_NSPoint=ff}fffI@{_NSSize=ff}{?=b1b1b1}}4@4:8 */
struct _NSTypesetterGlyphInfo {
	struct _NSPoint field_0;
	float field_1;
	float field_2;
	float field_3;
	unsigned int field_4;
	id field_5;
	struct _NSSize field_6;
	struct pyobjcanonymous0 field_7;
};

static struct _NSTypesetterGlyphInfo  *
meth_imp_355(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSTypesetterGlyphInfo  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSTypesetterGlyphInfo={_NSPoint=ff}fffI@{_NSSize=ff}{pyobjcanonymous0=ss}}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_355(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSTypesetterGlyphInfo  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct _NSTypesetterGlyphInfo  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSTypesetterGlyphInfo={_NSPoint=ff}fffI@{_NSSize=ff}{pyobjcanonymous0=ss}}", &objc_retval);
	return v;
}


/* signature: ^{_NSTypesetterGlyphInfo={_NSPoint=ff}fffI@{_NSSize=ff}{?=b1b1b1}}8@4:8i12 */
static struct _NSTypesetterGlyphInfo  *
meth_imp_356(id self, SEL sel, int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSTypesetterGlyphInfo  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSTypesetterGlyphInfo={_NSPoint=ff}fffI@{_NSSize=ff}{pyobjcanonymous0=ss}}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_356(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSTypesetterGlyphInfo  *objc_retval;
	int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _NSTypesetterGlyphInfo  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSTypesetterGlyphInfo={_NSPoint=ff}fffI@{_NSSize=ff}{pyobjcanonymous0=ss}}", &objc_retval);
	return v;
}


/* signature: ^{_NSZone=}4@4:8 */
struct _NSZone;
static struct _NSZone  *
meth_imp_357(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NSZone  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NSZone=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_357(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSZone  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct _NSZone  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NSZone=}", &objc_retval);
	return v;
}


/* signature: ^{_NXStream=I**iilii^{stream_functions}^v}4@4:8 */
struct _NXStream;
static struct _NXStream  *
meth_imp_358(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _NXStream  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_NXStream=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_358(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NXStream  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct _NXStream  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_NXStream=}", &objc_retval);
	return v;
}


/* signature: ^{_PrivatePrintOperationInfo={_NSRect={_NSPoint=ff}{_NSSize=ff}}{_NSRect={_NSPoint=ff}{_NSSize=ff}}cccccccciiiiiii@@{_NSRect={_NSPoint=ff}{_NSSize=ff}}ccciffffii{_NSPoint=ff}I^{_NSModalSession}@iiciii@c@ic@@i@}4@4:8 */
struct _NSModalSession;struct _PrivatePrintOperationInfo {
	struct _NSRect field_0;
	struct _NSRect field_1;
	char field_2;
	char field_3;
	char field_4;
	char field_5;
	char field_6;
	char field_7;
	char field_8;
	char field_9;
	int field_10;
	int field_11;
	int field_12;
	int field_13;
	int field_14;
	int field_15;
	int field_16;
	id field_17;
	id field_18;
	struct _NSRect field_19;
	char field_20;
	char field_21;
	char field_22;
	int field_23;
	float field_24;
	float field_25;
	float field_26;
	float field_27;
	int field_28;
	int field_29;
	struct _NSPoint field_30;
	unsigned int field_31;
	struct _NSModalSession  *field_32;
	id field_33;
	int field_34;
	int field_35;
	char field_36;
	int field_37;
	int field_38;
	int field_39;
	id field_40;
	char field_41;
	id field_42;
	int field_43;
	char field_44;
	id field_45;
	id field_46;
	int field_47;
	id field_48;
};

static struct _PrivatePrintOperationInfo  *
meth_imp_359(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _PrivatePrintOperationInfo  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_PrivatePrintOperationInfo={_NSRect={_NSPoint=ff}{_NSSize=ff}}{_NSRect={_NSPoint=ff}{_NSSize=ff}}cccccccciiiiiii@@{_NSRect={_NSPoint=ff}{_NSSize=ff}}ccciffffii{_NSPoint=ff}I^{_NSModalSession=}@iiciii@c@ic@@i@}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_359(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _PrivatePrintOperationInfo  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct _PrivatePrintOperationInfo  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_PrivatePrintOperationInfo={_NSRect={_NSPoint=ff}{_NSSize=ff}}{_NSRect={_NSPoint=ff}{_NSSize=ff}}cccccccciiiiiii@@{_NSRect={_NSPoint=ff}{_NSSize=ff}}ccciffffii{_NSPoint=ff}I^{_NSModalSession=}@iiciii@c@ic@@i@}", &objc_retval);
	return v;
}


/* signature: ^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}12@4:8^{OpaqueIconRef=}12i16 */
struct _RepresentationInfo;
struct OpaqueIconRef;
static struct _RepresentationInfo  *
meth_imp_360(id self, SEL sel, struct OpaqueIconRef  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _RepresentationInfo  *objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{OpaqueIconRef=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_RepresentationInfo=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_360(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _RepresentationInfo  *objc_retval;
	struct OpaqueIconRef  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{OpaqueIconRef=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _RepresentationInfo  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_RepresentationInfo=}", &objc_retval);
	return v;
}


/* signature: ^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}16@4:8i12@16@20 */
struct _RepresentationInfo;
static struct _RepresentationInfo  *
meth_imp_361(id self, SEL sel, int arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _RepresentationInfo  *objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_RepresentationInfo=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_361(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _RepresentationInfo  *objc_retval;
	int objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _RepresentationInfo  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_RepresentationInfo=}", &objc_retval);
	return v;
}


/* signature: ^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}32@4:8c12@16f36c24 */
struct _RepresentationInfo;
static struct _RepresentationInfo  *
meth_imp_362(id self, SEL sel, char arg_2, id arg_3, float arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _RepresentationInfo  *objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_RepresentationInfo=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_362(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _RepresentationInfo  *objc_retval;
	char objc_arg2;
	id objc_arg3;
	float objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _RepresentationInfo  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_RepresentationInfo=}", &objc_retval);
	return v;
}


/* signature: ^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}8@4:8@12 */
struct _RepresentationInfo;
static struct _RepresentationInfo  *
meth_imp_363(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _RepresentationInfo  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_RepresentationInfo=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_363(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _RepresentationInfo  *objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _RepresentationInfo  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_RepresentationInfo=}", &objc_retval);
	return v;
}


/* signature: ^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}12@4:8i12^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}16 */
struct _RowEntry;
struct _RowEntry;
static struct _RowEntry  *
meth_imp_364(id self, SEL sel, int arg_2, struct _RowEntry  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _RowEntry  *objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_RowEntry=}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_RowEntry=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_364(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _RowEntry  *objc_retval;
	int objc_arg2;
	struct _RowEntry  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_RowEntry=}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _RowEntry  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_RowEntry=}", &objc_retval);
	return v;
}


/* signature: ^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}13@4:8^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}12@16c20 */
struct _RowEntry;
struct _RowEntry;
static struct _RowEntry  *
meth_imp_365(id self, SEL sel, struct _RowEntry  *arg_2, id arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _RowEntry  *objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_RowEntry=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_RowEntry=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_365(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _RowEntry  *objc_retval;
	struct _RowEntry  *objc_arg2;
	id objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_RowEntry=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _RowEntry  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_RowEntry=}", &objc_retval);
	return v;
}


/* signature: ^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}20@4:8^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}12c16c20i24 */
struct _RowEntry;
struct _RowEntry;
static struct _RowEntry  *
meth_imp_366(id self, SEL sel, struct _RowEntry  *arg_2, char arg_3, char arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _RowEntry  *objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_RowEntry=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_RowEntry=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_366(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _RowEntry  *objc_retval;
	struct _RowEntry  *objc_arg2;
	char objc_arg3;
	char objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_RowEntry=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _RowEntry  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_RowEntry=}", &objc_retval);
	return v;
}


/* signature: ^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}8@4:8@12 */
struct _RowEntry;
static struct _RowEntry  *
meth_imp_367(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _RowEntry  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_RowEntry=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_367(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _RowEntry  *objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _RowEntry  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_RowEntry=}", &objc_retval);
	return v;
}


/* signature: ^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}8@4:8i12 */
struct _RowEntry;
static struct _RowEntry  *
meth_imp_368(id self, SEL sel, int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct _RowEntry  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{_RowEntry=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_368(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _RowEntry  *objc_retval;
	int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct _RowEntry  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{_RowEntry=}", &objc_retval);
	return v;
}


/* signature: ^{__CFArray=}5@4:8c12 */
struct __CFArray;
static struct __CFArray  *
meth_imp_369(id self, SEL sel, char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct __CFArray  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{__CFArray=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_369(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFArray  *objc_retval;
	char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct __CFArray  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{__CFArray=}", &objc_retval);
	return v;
}


/* signature: ^{__CFArray=}8@4:8@12 */
struct __CFArray;
static struct __CFArray  *
meth_imp_370(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct __CFArray  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{__CFArray=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_370(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFArray  *objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct __CFArray  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{__CFArray=}", &objc_retval);
	return v;
}


/* signature: ^{__CFDate=}4@4:8 */
struct __CFDate;
static struct __CFDate  *
meth_imp_371(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct __CFDate  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{__CFDate=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_371(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFDate  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct __CFDate  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{__CFDate=}", &objc_retval);
	return v;
}


/* signature: ^{__CFDictionary=}8@4:8@12 */
struct __CFDictionary;
static struct __CFDictionary  *
meth_imp_372(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct __CFDictionary  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{__CFDictionary=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_372(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFDictionary  *objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct __CFDictionary  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{__CFDictionary=}", &objc_retval);
	return v;
}


/* signature: ^{__CFHTTPMessage=}9@4:8@12c16 */
struct __CFHTTPMessage;
static struct __CFHTTPMessage  *
meth_imp_373(id self, SEL sel, id arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct __CFHTTPMessage  *objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{__CFHTTPMessage=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_373(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFHTTPMessage  *objc_retval;
	id objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct __CFHTTPMessage  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{__CFHTTPMessage=}", &objc_retval);
	return v;
}


/* signature: ^{__CFNotificationCenter=}4@4:8 */
struct __CFNotificationCenter;
static struct __CFNotificationCenter  *
meth_imp_374(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct __CFNotificationCenter  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{__CFNotificationCenter=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_374(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFNotificationCenter  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct __CFNotificationCenter  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{__CFNotificationCenter=}", &objc_retval);
	return v;
}


/* signature: ^{__CFPasteboard=}4@4:8 */
struct __CFPasteboard;
static struct __CFPasteboard  *
meth_imp_375(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct __CFPasteboard  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{__CFPasteboard=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_375(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFPasteboard  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct __CFPasteboard  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{__CFPasteboard=}", &objc_retval);
	return v;
}


/* signature: ^{__CFRunLoop=}4@4:8 */
struct __CFRunLoop;
static struct __CFRunLoop  *
meth_imp_376(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct __CFRunLoop  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{__CFRunLoop=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_376(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFRunLoop  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct __CFRunLoop  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{__CFRunLoop=}", &objc_retval);
	return v;
}


/* signature: ^{__CFSet=}5@4:8c12 */
struct __CFSet;
static struct __CFSet  *
meth_imp_377(id self, SEL sel, char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct __CFSet  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{__CFSet=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_377(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFSet  *objc_retval;
	char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct __CFSet  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{__CFSet=}", &objc_retval);
	return v;
}


/* signature: ^{__CFSocket=}8@4:8@12 */
struct __CFSocket;
static struct __CFSocket  *
meth_imp_378(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct __CFSocket  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{__CFSocket=}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_378(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFSocket  *objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct __CFSocket  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{__CFSocket=}", &objc_retval);
	return v;
}


/* signature: ^{__EventHandlerInfo=@:}12@4:8I12I16 */
struct __EventHandlerInfo {
	id field_0;
	SEL field_1;
};

static struct __EventHandlerInfo  *
meth_imp_379(id self, SEL sel, unsigned int arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct __EventHandlerInfo  *objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{__EventHandlerInfo=@:}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_379(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __EventHandlerInfo  *objc_retval;
	unsigned int objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct __EventHandlerInfo  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{__EventHandlerInfo=@:}", &objc_retval);
	return v;
}


/* signature: ^{objc_method_description=:*}8@4:8:12 */
struct objc_method_description {
	SEL field_0;
	char* field_1;
};

static struct objc_method_description  *
meth_imp_380(id self, SEL sel, SEL arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct objc_method_description  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{objc_method_description=:*}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_380(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct objc_method_description  *objc_retval;
	SEL objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (struct objc_method_description  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{objc_method_description=:*}", &objc_retval);
	return v;
}


/* signature: c12@4:8#12@16 */
static char 
meth_imp_381(id self, SEL sel, Class arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_381(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	Class objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8*12I16 */
static char 
meth_imp_382(id self, SEL sel, char* arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_382(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	char* objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8:12@16 */
static char 
meth_imp_383(id self, SEL sel, SEL arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_383(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	SEL objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8@12:16 */
static char 
meth_imp_384(id self, SEL sel, id arg_2, SEL arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_384(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	SEL objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8@12@16 */
static char 
meth_imp_385(id self, SEL sel, id arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_385(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8@12I16 */
static char 
meth_imp_386(id self, SEL sel, id arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_386(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8@12^@16 */
static char 
meth_imp_387(id self, SEL sel, id arg_2, id  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_387(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8@12^c16 */
static char 
meth_imp_388(id self, SEL sel, id arg_2, char  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_388(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	char  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8@12^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}16 */
struct _RepresentationInfo;
static char 
meth_imp_389(id self, SEL sel, id arg_2, struct _RepresentationInfo  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_RepresentationInfo=}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_389(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _RepresentationInfo  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_RepresentationInfo=}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8@12i16 */
static char 
meth_imp_390(id self, SEL sel, id arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_390(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8@12r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
static char 
meth_imp_391(id self, SEL sel, id arg_2, struct _NSRect  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_391(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSRect  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8I12I16 */
static char 
meth_imp_392(id self, SEL sel, unsigned int arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_392(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	unsigned int objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8^@12@16 */
static char 
meth_imp_393(id self, SEL sel, id  *arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_393(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id  *objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8^@12I16 */
static char 
meth_imp_394(id self, SEL sel, id  *arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_394(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id  *objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8^@12^I16 */
static char 
meth_imp_395(id self, SEL sel, id  *arg_2, unsigned int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_395(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id  *objc_arg2;
	unsigned int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8^{FSRef=[80C]}12@16 */
static char 
meth_imp_396(id self, SEL sel, struct FSRef  *arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_396(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct FSRef  *objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8^{tiff=*^{_NXStream}sccsll{?=IIIIIISSSSSSSSSSIIIffSSffII[2S]ISSSSI^S^S^S^S[3^S]*********[2I]II^I^I[2S]^f[2S]S^f^f^f[4^S]S[2S]**I^v}{?=SSL}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}12i16 */
static char 
meth_imp_397(id self, SEL sel, struct tiff  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{tiff=*^{_NXStream=}sccsll{pyobjcanonymous0=ss}{pyobjcanonymous0=ss}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_397(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct tiff  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{tiff=*^{_NXStream=}sccsll{pyobjcanonymous0=ss}{pyobjcanonymous0=ss}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8i12@16 */
static char 
meth_imp_398(id self, SEL sel, int arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_398(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8i12i16 */
static char 
meth_imp_399(id self, SEL sel, int arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_399(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@16 */
static char 
meth_imp_400(id self, SEL sel, struct _NSRect  *arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_400(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSRect  *objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8{NSButtonState=iccc}12 */
static char 
meth_imp_401(id self, SEL sel, struct NSButtonState arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{NSButtonState=iccc}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_401(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct NSButtonState objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{NSButtonState=iccc}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c12@4:8{_NSPoint=ff}12 */
static char 
meth_imp_402(id self, SEL sel, struct _NSPoint arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_402(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSPoint objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c13@4:8@12@16c20 */
static char 
meth_imp_403(id self, SEL sel, id arg_2, id arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_403(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c13@4:8@12c16c20 */
static char 
meth_imp_404(id self, SEL sel, id arg_2, char arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_404(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	char objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c14@4:8@12@16S20 */
static char 
meth_imp_405(id self, SEL sel, id arg_2, id arg_3, unsigned short arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_405(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	unsigned short objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8*12I16@20 */
static char 
meth_imp_406(id self, SEL sel, char* arg_2, unsigned int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_406(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	char* objc_arg2;
	unsigned int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8*12I16I20 */
static char 
meth_imp_407(id self, SEL sel, char* arg_2, unsigned int arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_407(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	char* objc_arg2;
	unsigned int objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8:12@16@20 */
static char 
meth_imp_408(id self, SEL sel, SEL arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_408(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	SEL objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12@16:20 */
static char 
meth_imp_409(id self, SEL sel, id arg_2, id arg_3, SEL arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_409(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	SEL objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12@16@20 */
static char 
meth_imp_410(id self, SEL sel, id arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_410(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12@16I20 */
static char 
meth_imp_411(id self, SEL sel, id arg_2, id arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_411(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12@16^c20 */
static char 
meth_imp_412(id self, SEL sel, id arg_2, id arg_3, char  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_412(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	char  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12@16i20 */
static char 
meth_imp_413(id self, SEL sel, id arg_2, id arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_413(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12^@16^@20 */
static char 
meth_imp_414(id self, SEL sel, id arg_2, id  *arg_3, id  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_414(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id  *objc_arg3;
	id  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16^c20 */
static char 
meth_imp_415(id self, SEL sel, id arg_2, struct _NSRect  *arg_3, char  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_415(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSRect  *objc_arg3;
	char  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12i16i20 */
static char 
meth_imp_416(id self, SEL sel, id arg_2, int arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_416(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	int objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12r^{FSRef=[80C]}16r^{FSRef=[80C]}20 */
static char 
meth_imp_417(id self, SEL sel, id arg_2, struct FSRef  *arg_3, struct FSRef  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_417(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct FSRef  *objc_arg3;
	struct FSRef  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16i20 */
static char 
meth_imp_418(id self, SEL sel, id arg_2, struct _NSRect  *arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_418(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSRect  *objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12{_NSPoint=ff}16 */
static char 
meth_imp_419(id self, SEL sel, id arg_2, struct _NSPoint arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_419(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSPoint objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8@12{_NSRange=II}16 */
static char 
meth_imp_420(id self, SEL sel, id arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_420(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8I12I16@20 */
static char 
meth_imp_421(id self, SEL sel, unsigned int arg_2, unsigned int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_421(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	unsigned int objc_arg2;
	unsigned int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8^@12@16^@20 */
static char 
meth_imp_422(id self, SEL sel, id  *arg_2, id arg_3, id  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_422(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id  *objc_arg2;
	id objc_arg3;
	id  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8^I12^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@20 */
static char 
meth_imp_423(id self, SEL sel, unsigned int  *arg_2, struct _NSRect  *arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_423(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	unsigned int  *objc_arg2;
	struct _NSRect  *objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8^i12^i16@20 */
static char 
meth_imp_424(id self, SEL sel, int  *arg_2, int  *arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_424(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int  *objc_arg2;
	int  *objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8i12@16@20 */
static char 
meth_imp_425(id self, SEL sel, int arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_425(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8i12i16i20 */
static char 
meth_imp_426(id self, SEL sel, int arg_2, int arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_426(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int objc_arg2;
	int objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8s12r^{FSRef=[80C]}16^{FSRef=[80C]}20 */
static char 
meth_imp_427(id self, SEL sel, short arg_2, struct FSRef  *arg_3, struct FSRef  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_427(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	short objc_arg2;
	struct FSRef  *objc_arg3;
	struct FSRef  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8{_NSPoint=ff}12@20 */
static char 
meth_imp_428(id self, SEL sel, struct _NSPoint arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_428(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSPoint objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c16@4:8{_NSPoint=ff}12i20 */
static char 
meth_imp_429(id self, SEL sel, struct _NSPoint arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_429(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSPoint objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c17@4:8@12^{FSRef=[80C]}16c20c24 */
static char 
meth_imp_430(id self, SEL sel, id arg_2, struct FSRef  *arg_3, char arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_430(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct FSRef  *objc_arg3;
	char objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c20@4:8:12@16i20i24 */
static char 
meth_imp_431(id self, SEL sel, SEL arg_2, id arg_3, int arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_431(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	SEL objc_arg2;
	id objc_arg3;
	int objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c20@4:8@12@16@20I24 */
static char 
meth_imp_432(id self, SEL sel, id arg_2, id arg_3, id arg_4, unsigned int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_432(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	unsigned int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c20@4:8@12@16@20i24 */
static char 
meth_imp_433(id self, SEL sel, id arg_2, id arg_3, id arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_433(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c20@4:8@12{_NSRange=II}16@24 */
static char 
meth_imp_434(id self, SEL sel, id arg_2, struct _NSRange arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_434(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSRange objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c20@4:8^@12@16I20@24 */
static char 
meth_imp_435(id self, SEL sel, id  *arg_2, id arg_3, unsigned int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_435(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id  *objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c20@4:8^i12^i16@20r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}24 */
static char 
meth_imp_436(id self, SEL sel, int  *arg_2, int  *arg_3, id arg_4, struct _NSRect  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_436(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int  *objc_arg2;
	int  *objc_arg3;
	id objc_arg4;
	struct _NSRect  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c20@4:8^i12^i16{_NSPoint=ff}20 */
static char 
meth_imp_437(id self, SEL sel, int  *arg_2, int  *arg_3, struct _NSPoint arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_437(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int  *objc_arg2;
	int  *objc_arg3;
	struct _NSPoint objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c20@4:8i12@16@20@24 */
static char 
meth_imp_438(id self, SEL sel, int arg_2, id arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_438(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c20@4:8{_NSPoint=ff}12^i20^i24 */
static char 
meth_imp_439(id self, SEL sel, struct _NSPoint arg_2, int  *arg_3, int  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_439(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSPoint objc_arg2;
	int  *objc_arg3;
	int  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12 */
static char 
meth_imp_440(id self, SEL sel, struct _NSRect arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_440(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSRect objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c21@4:8*12i16c20c24c28 */
static char 
meth_imp_441(id self, SEL sel, char* arg_2, int arg_3, char arg_4, char arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_441(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	char* objc_arg2;
	int objc_arg3;
	char objc_arg4;
	char objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c21@4:8@12@16c20c24c28 */
static char 
meth_imp_442(id self, SEL sel, id arg_2, id arg_3, char arg_4, char arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_442(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	char objc_arg4;
	char objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c21@4:8@12I16^@20@24c28 */
static char 
meth_imp_443(id self, SEL sel, id arg_2, unsigned int arg_3, id  *arg_4, id arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_443(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	id  *objc_arg4;
	id objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c24@4:8@12@16@20@24^i28 */
static char 
meth_imp_444(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, int  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_444(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	int  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c24@4:8@12@16i20^{_NSMapTable=}24@28 */
struct _NSMapTable;
static char 
meth_imp_445(id self, SEL sel, id arg_2, id arg_3, int arg_4, struct _NSMapTable  *arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSMapTable=}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_445(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	struct _NSMapTable  *objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSMapTable=}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c24@4:8@12@16{_NSPoint=ff}20@28 */
static char 
meth_imp_446(id self, SEL sel, id arg_2, id arg_3, struct _NSPoint arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_446(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct _NSPoint objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c24@4:8@12I16@20@24I28 */
static char 
meth_imp_447(id self, SEL sel, id arg_2, unsigned int arg_3, id arg_4, id arg_5, unsigned int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_447(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	id objc_arg4;
	id objc_arg5;
	unsigned int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c24@4:8@12i16^c20^c24^@28 */
static char 
meth_imp_448(id self, SEL sel, id arg_2, int arg_3, char  *arg_4, char  *arg_5, id  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_448(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	int objc_arg3;
	char  *objc_arg4;
	char  *objc_arg5;
	id  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c24@4:8@12r^{FSRef=[80C]}16r^{FSRef=[80C]}20@24i28 */
static char 
meth_imp_449(id self, SEL sel, id arg_2, struct FSRef  *arg_3, struct FSRef  *arg_4, id arg_5, int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_449(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct FSRef  *objc_arg3;
	struct FSRef  *objc_arg4;
	id objc_arg5;
	int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c24@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
static char 
meth_imp_450(id self, SEL sel, id arg_2, struct _NSRect arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_450(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSRect objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c24@4:8I12{_NSPoint=ff}16I24@28 */
static char 
meth_imp_451(id self, SEL sel, unsigned int arg_2, struct _NSPoint arg_3, unsigned int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_451(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	unsigned int objc_arg2;
	struct _NSPoint objc_arg3;
	unsigned int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c24@4:8{_NSPoint=ff}12{_NSPoint=ff}20@28 */
static char 
meth_imp_452(id self, SEL sel, struct _NSPoint arg_2, struct _NSPoint arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_452(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSPoint objc_arg2;
	struct _NSPoint objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c24@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28 */
static char 
meth_imp_453(id self, SEL sel, struct _NSRect arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_453(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSRect objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c25@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16c32 */
static char 
meth_imp_454(id self, SEL sel, id arg_2, struct _NSRect arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_454(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSRect objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c25@4:8^i12@16@20i24c28c32 */
static char 
meth_imp_455(id self, SEL sel, int  *arg_2, id arg_3, id arg_4, int arg_5, char arg_6, char arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_455(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int  *objc_arg2;
	id objc_arg3;
	id objc_arg4;
	int objc_arg5;
	char objc_arg6;
	char objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c28@4:8@12^c16^c20^c24^@28^@32 */
static char 
meth_imp_456(id self, SEL sel, id arg_2, char  *arg_3, char  *arg_4, char  *arg_5, id  *arg_6, id  *arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_456(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	char  *objc_arg3;
	char  *objc_arg4;
	char  *objc_arg5;
	id  *objc_arg6;
	id  *objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c28@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32 */
static char 
meth_imp_457(id self, SEL sel, id arg_2, struct _NSRect arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_457(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c28@4:8^@12^{_NSRange=II}16@20{_NSRange=II}24^@32 */
static char 
meth_imp_458(id self, SEL sel, id  *arg_2, struct _NSRange  *arg_3, id arg_4, struct _NSRange arg_5, id  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_458(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id  *objc_arg2;
	struct _NSRange  *objc_arg3;
	id objc_arg4;
	struct _NSRange objc_arg5;
	id  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c28@4:8{_NSPoint=ff}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}20 */
static char 
meth_imp_459(id self, SEL sel, struct _NSPoint arg_2, struct _NSRect arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_459(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSPoint objc_arg2;
	struct _NSRect objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32 */
static char 
meth_imp_460(id self, SEL sel, struct _NSRect arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_460(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSRect objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c32@4:8^i12{_NSSize=ff}16f36 */
static char 
meth_imp_461(id self, SEL sel, int  *arg_2, struct _NSSize arg_3, float arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_461(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int  *objc_arg2;
	struct _NSSize objc_arg3;
	float objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c32@4:8f36 */
static char 
meth_imp_462(id self, SEL sel, float arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_462(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	float objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c32@4:8f36c16 */
static char 
meth_imp_463(id self, SEL sel, float arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_463(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	float objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c32@4:8i12f36r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}20r^{_NSPoint=ff}24 */
static char 
meth_imp_464(id self, SEL sel, int arg_2, float arg_3, struct _NSRect  *arg_4, struct _NSPoint  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_464(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int objc_arg2;
	float objc_arg3;
	struct _NSRect  *objc_arg4;
	struct _NSPoint  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c32@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12f36 */
static char 
meth_imp_465(id self, SEL sel, struct _NSRect  *arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_465(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSRect  *objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c36@4:8@12^{FSRef=[80C]}16@20^{FSRef=[80C]}24i28^{_NSMapTable=}32@40 */
struct _NSMapTable;
static char 
meth_imp_466(id self, SEL sel, id arg_2, struct FSRef  *arg_3, id arg_4, struct FSRef  *arg_5, int arg_6, struct _NSMapTable  *arg_7, id arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("^{_NSMapTable=}", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_466(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct FSRef  *objc_arg3;
	id objc_arg4;
	struct FSRef  *objc_arg5;
	int objc_arg6;
	struct _NSMapTable  *objc_arg7;
	id objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("^{_NSMapTable=}", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c36@4:8@12i16i20c24c28c32c43 */
static char 
meth_imp_467(id self, SEL sel, id arg_2, int arg_3, int arg_4, char arg_5, char arg_6, char arg_7, char arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_467(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	int objc_arg3;
	int objc_arg4;
	char objc_arg5;
	char objc_arg6;
	char objc_arg7;
	char objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c36@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32I40 */
static char 
meth_imp_468(id self, SEL sel, id arg_2, struct _NSRect arg_3, id arg_4, unsigned int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_468(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	unsigned int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c36@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32c43 */
static char 
meth_imp_469(id self, SEL sel, id arg_2, struct _NSRect arg_3, id arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_469(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c36@4:8d36 */
static char 
meth_imp_470(id self, SEL sel, double arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_470(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	double objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c36@4:8d36^v20@24@28I32 */
static char 
meth_imp_471(id self, SEL sel, double arg_2, void  *arg_3, id arg_4, id arg_5, unsigned int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_471(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	double objc_arg2;
	void  *objc_arg3;
	id objc_arg4;
	id objc_arg5;
	unsigned int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c36@4:8{_NSRange=II}12{_NSRange=II}20{_NSRange=II}28@40 */
static char 
meth_imp_472(id self, SEL sel, struct _NSRange arg_2, struct _NSRange arg_3, struct _NSRange arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_472(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSRange objc_arg2;
	struct _NSRange objc_arg3;
	struct _NSRange objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28i32i40 */
static char 
meth_imp_473(id self, SEL sel, struct _NSRect arg_2, id arg_3, int arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_473(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSRect objc_arg2;
	id objc_arg3;
	int objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c40@4:8*12I16^I20I24c28{_NSRange=II}36^{_NSRange=II}44 */
static char 
meth_imp_474(id self, SEL sel, char* arg_2, unsigned int arg_3, unsigned int  *arg_4, unsigned int arg_5, char arg_6, struct _NSRange arg_7, struct _NSRange  *arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_474(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	char* objc_arg2;
	unsigned int objc_arg3;
	unsigned int  *objc_arg4;
	unsigned int objc_arg5;
	char objc_arg6;
	struct _NSRange objc_arg7;
	struct _NSRange  *objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c40@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32I40c47 */
static char 
meth_imp_475(id self, SEL sel, id arg_2, struct _NSRect arg_3, id arg_4, unsigned int arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_475(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	unsigned int objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c40@4:8^@12I16^I20I24c28{_NSRange=II}36^{_NSRange=II}44 */
static char 
meth_imp_476(id self, SEL sel, id  *arg_2, unsigned int arg_3, unsigned int  *arg_4, unsigned int arg_5, char arg_6, struct _NSRange arg_7, struct _NSRange  *arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_476(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id  *objc_arg2;
	unsigned int objc_arg3;
	unsigned int  *objc_arg4;
	unsigned int objc_arg5;
	char objc_arg6;
	struct _NSRange objc_arg7;
	struct _NSRange  *objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c40@4:8d36@20@24@28@32I40I44 */
static char 
meth_imp_477(id self, SEL sel, double arg_2, id arg_3, id arg_4, id arg_5, id arg_6, unsigned int arg_7, unsigned int arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_477(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	double objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	unsigned int objc_arg7;
	unsigned int objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c4@4:8 */
static char 
meth_imp_478(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_478(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c56@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32i48f36c59c63 */
static char 
meth_imp_479(id self, SEL sel, struct _NSRect arg_2, struct _NSRect arg_3, int arg_4, float arg_5, char arg_6, char arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_479(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSRect objc_arg2;
	struct _NSRect objc_arg3;
	int objc_arg4;
	float objc_arg5;
	char objc_arg6;
	char objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c5@4:8c12 */
static char 
meth_imp_480(id self, SEL sel, char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_480(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c6@4:8S12 */
static char 
meth_imp_481(id self, SEL sel, unsigned short arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_481(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	unsigned short objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c6@4:8s12 */
static char 
meth_imp_482(id self, SEL sel, short arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_482(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	short objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8#12 */
static char 
meth_imp_483(id self, SEL sel, Class arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_483(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	Class objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8:12 */
static char 
meth_imp_484(id self, SEL sel, SEL arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_484(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	SEL objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8@12 */
static char 
meth_imp_485(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_485(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8I12 */
static char 
meth_imp_486(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_486(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8L12 */
static char 
meth_imp_487(id self, SEL sel, unsigned long arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("L", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_487(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	unsigned long objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("L", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8^*12 */
static char 
meth_imp_488(id self, SEL sel, char*  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_488(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	char*  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8^I12 */
static char 
meth_imp_489(id self, SEL sel, unsigned int  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_489(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	unsigned int  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8^d12 */
static char 
meth_imp_490(id self, SEL sel, double  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_490(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	double  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8^f12 */
static char 
meth_imp_491(id self, SEL sel, float  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_491(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	float  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8^i12 */
static char 
meth_imp_492(id self, SEL sel, int  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_492(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8^q12 */
static char 
meth_imp_493(id self, SEL sel, long long  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^q", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_493(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	long long  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^q", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8^v12 */
static char 
meth_imp_494(id self, SEL sel, void  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_494(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	void  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8^{_NSPoint=ff}12 */
static char 
meth_imp_495(id self, SEL sel, struct _NSPoint  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_495(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSPoint  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}12 */
struct _RepresentationInfo;
static char 
meth_imp_496(id self, SEL sel, struct _RepresentationInfo  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_RepresentationInfo=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_496(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _RepresentationInfo  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_RepresentationInfo=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8i12 */
static char 
meth_imp_497(id self, SEL sel, int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_497(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8r*12 */
static char 
meth_imp_498(id self, SEL sel, char* arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_498(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	char* objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8r^{FSRef=[80C]}12 */
static char 
meth_imp_499(id self, SEL sel, struct FSRef  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_499(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct FSRef  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c8@4:8r^{_NSPoint=ff}12 */
static char 
meth_imp_500(id self, SEL sel, struct _NSPoint  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_500(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSPoint  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c9@4:8@12c16 */
static char 
meth_imp_501(id self, SEL sel, id arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_501(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	id objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c9@4:8^{_NSPoint=ff}12c16 */
static char 
meth_imp_502(id self, SEL sel, struct _NSPoint  *arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_502(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSPoint  *objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c9@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c16 */
static char 
meth_imp_503(id self, SEL sel, struct _NSRect  *arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_503(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSRect  *objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c9@4:8^{_NSSize=ff}12c16 */
static char 
meth_imp_504(id self, SEL sel, struct _NSSize  *arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_504(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _NSSize  *objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c9@4:8^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}12c16 */
struct _RepresentationInfo;
static char 
meth_imp_505(id self, SEL sel, struct _RepresentationInfo  *arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_RepresentationInfo=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_505(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	struct _RepresentationInfo  *objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_RepresentationInfo=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: c9@4:8i12c16 */
static char 
meth_imp_506(id self, SEL sel, int arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("c", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_506(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_retval;
	int objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("c", &objc_retval);
	return v;
}


/* signature: d20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12 */
static double 
meth_imp_507(id self, SEL sel, struct _NSRect arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	double objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("d", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_507(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	double objc_retval;
	struct _NSRect objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (double)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("d", &objc_retval);
	return v;
}


/* signature: d36@4:8d36 */
static double 
meth_imp_508(id self, SEL sel, double arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	double objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("d", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_508(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	double objc_retval;
	double objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (double)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("d", &objc_retval);
	return v;
}


/* signature: d4@4:8 */
static double 
meth_imp_509(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	double objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("d", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_509(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	double objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (double)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("d", &objc_retval);
	return v;
}


/* signature: d8@4:8@12 */
static double 
meth_imp_510(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	double objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("d", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_510(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	double objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (double)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("d", &objc_retval);
	return v;
}


/* signature: d8@4:8i12 */
static double 
meth_imp_511(id self, SEL sel, int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	double objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("d", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_511(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	double objc_retval;
	int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (double)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("d", &objc_retval);
	return v;
}


/* signature: f12@4:8@12@16 */
static float 
meth_imp_512(id self, SEL sel, id arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_512(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f12@4:8@12I16 */
static float 
meth_imp_513(id self, SEL sel, id arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_513(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f12@4:8r*12I16 */
static float 
meth_imp_514(id self, SEL sel, char* arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_514(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	char* objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f12@4:8{_NSSize=ff}12 */
static float 
meth_imp_515(id self, SEL sel, struct _NSSize arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_515(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	struct _NSSize objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f16@4:8{_NSPoint=ff}12@20 */
static float 
meth_imp_516(id self, SEL sel, struct _NSPoint arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_516(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	struct _NSPoint objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f32@4:8@12@16f36 */
static float 
meth_imp_517(id self, SEL sel, id arg_2, id arg_3, float arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_517(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	id objc_arg2;
	id objc_arg3;
	float objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f32@4:8c12f36 */
static float 
meth_imp_518(id self, SEL sel, char arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_518(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	char objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f32@4:8f36 */
static float 
meth_imp_519(id self, SEL sel, float arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_519(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	float objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f36@4:8d36 */
static float 
meth_imp_520(id self, SEL sel, double arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_520(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	double objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f4@4:8 */
static float 
meth_imp_521(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_521(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f8@4:8@12 */
static float 
meth_imp_522(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_522(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f8@4:8I12 */
static float 
meth_imp_523(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_523(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: f8@4:8i12 */
static float 
meth_imp_524(id self, SEL sel, int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_524(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_retval;
	int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("f", &objc_retval);
	return v;
}


/* signature: i12@4:8*12@16 */
static int 
meth_imp_525(id self, SEL sel, char* arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_525(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	char* objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8@12:16 */
static int 
meth_imp_526(id self, SEL sel, id arg_2, SEL arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_526(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	SEL objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8@12@16 */
static int 
meth_imp_527(id self, SEL sel, id arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_527(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8@12I16 */
static int 
meth_imp_528(id self, SEL sel, id arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_528(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8@12^i16 */
static int 
meth_imp_529(id self, SEL sel, id arg_2, int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_529(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8@12i16 */
static int 
meth_imp_530(id self, SEL sel, id arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_530(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8S12i16 */
static int 
meth_imp_531(id self, SEL sel, unsigned short arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_531(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	unsigned short objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12^f16 */
static int 
meth_imp_532(id self, SEL sel, struct _NSRect  *arg_2, float  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_532(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct _NSRect  *objc_arg2;
	float  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8^{__sFILE=*iiss{__sbuf=*i}i^v^?^?^?^?{__sbuf=*i}*i[3C][1C]{__sbuf=*i}iq}12i16 */
static int 
meth_imp_533(id self, SEL sel, struct __sFILE  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{__sFILE=*iiss{__sbuf=*i}i^v^?^?^?^?{__sbuf=*i}*i[3C][1C]{__sbuf=*i}iq}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_533(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct __sFILE  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{__sFILE=*iiss{__sbuf=*i}i^v^?^?^?^?{__sbuf=*i}*i[3C][1C]{__sbuf=*i}iq}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8i12@16 */
static int 
meth_imp_534(id self, SEL sel, int arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_534(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	int objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8i12I16 */
static int 
meth_imp_535(id self, SEL sel, int arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_535(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	int objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8i12^{_NSPoint=ff}16 */
static int 
meth_imp_536(id self, SEL sel, int arg_2, struct _NSPoint  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_536(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	int objc_arg2;
	struct _NSPoint  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8i12i16 */
static int 
meth_imp_537(id self, SEL sel, int arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_537(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	int objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8r*12^i16 */
static int 
meth_imp_538(id self, SEL sel, char* arg_2, int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_538(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	char* objc_arg2;
	int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8{NSButtonState=iccc}12 */
static int 
meth_imp_539(id self, SEL sel, struct NSButtonState arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{NSButtonState=iccc}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_539(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct NSButtonState objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{NSButtonState=iccc}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i12@4:8{_NSPoint=ff}12 */
static int 
meth_imp_540(id self, SEL sel, struct _NSPoint arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_540(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct _NSPoint objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i13@4:8@12@16c20 */
static int 
meth_imp_541(id self, SEL sel, id arg_2, id arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_541(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	id objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i13@4:8@12i16c20 */
static int 
meth_imp_542(id self, SEL sel, id arg_2, int arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_542(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	int objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i16@4:8@12@16@20 */
static int 
meth_imp_543(id self, SEL sel, id arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_543(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i16@4:8@12@16i20 */
static int 
meth_imp_544(id self, SEL sel, id arg_2, id arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_544(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i16@4:8@12c16@20 */
static int 
meth_imp_545(id self, SEL sel, id arg_2, char arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_545(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	char objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i16@4:8@12{_NSRange=II}16 */
static int 
meth_imp_546(id self, SEL sel, id arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_546(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i16@4:8^I12i16^{_NSPoint=ff}20 */
static int 
meth_imp_547(id self, SEL sel, unsigned int  *arg_2, int arg_3, struct _NSPoint  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_547(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	unsigned int  *objc_arg2;
	int objc_arg3;
	struct _NSPoint  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i16@4:8i12c16@20 */
static int 
meth_imp_548(id self, SEL sel, int arg_2, char arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_548(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	int objc_arg2;
	char objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i16@4:8i12i16@20 */
static int 
meth_imp_549(id self, SEL sel, int arg_2, int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_549(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	int objc_arg2;
	int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i16@4:8i12{_NSPoint=ff}16 */
static int 
meth_imp_550(id self, SEL sel, int arg_2, struct _NSPoint arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_550(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	int objc_arg2;
	struct _NSPoint objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i17@4:8@12@16@20c24 */
static int 
meth_imp_551(id self, SEL sel, id arg_2, id arg_3, id arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_551(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i20@4:8@12@16@20@24 */
static int 
meth_imp_552(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_552(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i20@4:8@12I16{_NSRange=II}20 */
static int 
meth_imp_553(id self, SEL sel, id arg_2, unsigned int arg_3, struct _NSRange arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_553(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	struct _NSRange objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i20@4:8@12^S16^i20^{_NSSortState=iIIII[4@]}24 */
struct _NSSortState {
	int field_0;
	unsigned int field_1;
	unsigned int field_2;
	unsigned int field_3;
	unsigned int field_4;
	id field_5[4];
};

static int 
meth_imp_554(id self, SEL sel, id arg_2, unsigned short  *arg_3, int  *arg_4, struct _NSSortState  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^S", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSSortState=iIIII[4@]}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_554(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	unsigned short  *objc_arg3;
	int  *objc_arg4;
	struct _NSSortState  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^S", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSSortState=iIIII[4@]}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i20@4:8^{OpaqueEventRef=}12{Point=ss}16s20I24 */
struct OpaqueEventRef;
struct Point {
	short field_0;
	short field_1;
};

static int 
meth_imp_555(id self, SEL sel, struct OpaqueEventRef  *arg_2, struct Point arg_3, short arg_4, unsigned int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{OpaqueEventRef=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{Point=ss}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_555(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct OpaqueEventRef  *objc_arg2;
	struct Point objc_arg3;
	short objc_arg4;
	unsigned int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{OpaqueEventRef=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{Point=ss}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i20@4:8c12@16@20@24 */
static int 
meth_imp_556(id self, SEL sel, char arg_2, id arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_556(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	char objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12 */
static int 
meth_imp_557(id self, SEL sel, struct _NSRect arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_557(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct _NSRect objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i24@4:8@12@16@20@24^@28 */
static int 
meth_imp_558(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, id  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_558(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i24@4:8@12I16{_NSRange=II}20@28 */
static int 
meth_imp_559(id self, SEL sel, id arg_2, unsigned int arg_3, struct _NSRange arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_559(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	unsigned int objc_arg3;
	struct _NSRange objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i24@4:8@12c16@20@24@28 */
static int 
meth_imp_560(id self, SEL sel, id arg_2, char arg_3, id arg_4, id arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_560(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	char objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i24@4:8i12{_NSPoint=ff}16@24i28 */
static int 
meth_imp_561(id self, SEL sel, int arg_2, struct _NSPoint arg_3, id arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_561(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	int objc_arg2;
	struct _NSPoint objc_arg3;
	id objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i28@4:8@12@16@20@24@28@32 */
static int 
meth_imp_562(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, id arg_6, id arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_562(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	id objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28^v32 */
static int 
meth_imp_563(id self, SEL sel, struct _NSRect arg_2, id arg_3, void  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_563(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct _NSRect objc_arg2;
	id objc_arg3;
	void  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i32@4:8f36 */
static int 
meth_imp_564(id self, SEL sel, float arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_564(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	float objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i32@4:8i12f36 */
static int 
meth_imp_565(id self, SEL sel, int arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_565(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	int objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i36@4:8@12@16i20c24c28c32c43 */
static int 
meth_imp_566(id self, SEL sel, id arg_2, id arg_3, int arg_4, char arg_5, char arg_6, char arg_7, char arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_566(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	char objc_arg5;
	char objc_arg6;
	char objc_arg7;
	char objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i36@4:8@12{_NSRange=II}16@24{_NSRange=II}28i40 */
static int 
meth_imp_567(id self, SEL sel, id arg_2, struct _NSRange arg_3, id arg_4, struct _NSRange arg_5, int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_567(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	struct _NSRange objc_arg3;
	id objc_arg4;
	struct _NSRange objc_arg5;
	int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i36@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32^v40 */
static int 
meth_imp_568(id self, SEL sel, id arg_2, struct _NSRect arg_3, id arg_4, void  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_568(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	void  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i36@4:8d36 */
static int 
meth_imp_569(id self, SEL sel, double arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_569(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	double objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28^v32c43 */
static int 
meth_imp_570(id self, SEL sel, struct _NSRect arg_2, id arg_3, void  *arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_570(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct _NSRect objc_arg2;
	id objc_arg3;
	void  *objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28@32^v40 */
static int 
meth_imp_571(id self, SEL sel, struct _NSRect arg_2, char arg_3, id arg_4, void  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_571(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct _NSRect objc_arg2;
	char objc_arg3;
	id objc_arg4;
	void  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28@32@40@44 */
static int 
meth_imp_572(id self, SEL sel, struct _NSRect arg_2, char arg_3, id arg_4, id arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_572(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct _NSRect objc_arg2;
	char objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i48@4:8@12@16@20{_NSRect={_NSPoint=ff}{_NSSize=ff}}28@44c51^v52 */
static int 
meth_imp_573(id self, SEL sel, id arg_2, id arg_3, id arg_4, struct _NSRect arg_5, id arg_6, char arg_7, void  *arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_573(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct _NSRect objc_arg5;
	id objc_arg6;
	char objc_arg7;
	void  *objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i4@4:8 */
static int 
meth_imp_574(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_574(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i5@4:8c12 */
static int 
meth_imp_575(id self, SEL sel, char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_575(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i6@4:8S12 */
static int 
meth_imp_576(id self, SEL sel, unsigned short arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_576(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	unsigned short objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i8@4:8*12 */
static int 
meth_imp_577(id self, SEL sel, char* arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_577(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	char* objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i8@4:8@12 */
static int 
meth_imp_578(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_578(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i8@4:8I12 */
static int 
meth_imp_579(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_579(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i8@4:8^@12 */
static int 
meth_imp_580(id self, SEL sel, id  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_580(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i8@4:8^I12 */
static int 
meth_imp_581(id self, SEL sel, unsigned int  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_581(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	unsigned int  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i8@4:8^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}12 */
struct _NSModalSession;
static int 
meth_imp_582(id self, SEL sel, struct _NSModalSession  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSModalSession=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_582(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct _NSModalSession  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSModalSession=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i8@4:8i12 */
static int 
meth_imp_583(id self, SEL sel, int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_583(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i8@4:8r^{_NSPoint=ff}12 */
static int 
meth_imp_584(id self, SEL sel, struct _NSPoint  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_584(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	struct _NSPoint  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: i9@4:8@12c16 */
static int 
meth_imp_585(id self, SEL sel, id arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_585(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_retval;
	id objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (int)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("i", &objc_retval);
	return v;
}


/* signature: l4@4:8 */
static long 
meth_imp_586(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	long objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("l", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_586(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	long objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (long)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("l", &objc_retval);
	return v;
}


/* signature: q4@4:8 */
static long long 
meth_imp_587(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	long long objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("q", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_587(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	long long objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (long long)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("q", &objc_retval);
	return v;
}


/* signature: q8@4:8@12 */
static long long 
meth_imp_588(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	long long objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("q", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_588(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	long long objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (long long)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("q", &objc_retval);
	return v;
}


/* signature: r*4@4:8 */
static char* 
meth_imp_589(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char* objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("*", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_589(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (char*)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("*", &objc_retval);
	return v;
}


/* signature: r*5@4:8c12 */
static char* 
meth_imp_590(id self, SEL sel, char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char* objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("*", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_590(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_retval;
	char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char*)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("*", &objc_retval);
	return v;
}


/* signature: r*8@4:8@12 */
static char* 
meth_imp_591(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char* objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("*", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_591(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char*)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("*", &objc_retval);
	return v;
}


/* signature: r*8@4:8I12 */
static char* 
meth_imp_592(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	char* objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("*", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_592(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_retval;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (char*)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("*", &objc_retval);
	return v;
}


/* signature: r^I4@4:8 */
static unsigned int  *
meth_imp_593(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	unsigned int  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^I", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_593(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (unsigned int  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^I", &objc_retval);
	return v;
}


/* signature: r^f4@4:8 */
static float  *
meth_imp_594(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_594(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (float  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^f", &objc_retval);
	return v;
}


/* signature: r^f8@4:8@12 */
static float  *
meth_imp_595(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	float  *objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^f", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_595(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float  *objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (float  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^f", &objc_retval);
	return v;
}


/* signature: r^i4@4:8 */
static int  *
meth_imp_596(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	int  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^i", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_596(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (int  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^i", &objc_retval);
	return v;
}


/* signature: r^v4@4:8 */
static void  *
meth_imp_597(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	void  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^v", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_597(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (void  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^v", &objc_retval);
	return v;
}


/* signature: r^{FSRef=[80C]}4@4:8 */
static struct FSRef  *
meth_imp_598(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	struct FSRef  *objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_598(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct FSRef  *objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (struct FSRef  *)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("^{FSRef=[80C]}", &objc_retval);
	return v;
}


/* signature: s12@4:8@12@16 */
static short 
meth_imp_599(id self, SEL sel, id arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	short objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("s", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_599(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	short objc_retval;
	id objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (short)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("s", &objc_retval);
	return v;
}


/* signature: s12@4:8L12@16 */
static short 
meth_imp_600(id self, SEL sel, unsigned long arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	short objc_retval;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("L", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("s", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_600(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	short objc_retval;
	unsigned long objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("L", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (short)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("s", &objc_retval);
	return v;
}


/* signature: s16@4:8@12@16@20 */
static short 
meth_imp_601(id self, SEL sel, id arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	short objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("s", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_601(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	short objc_retval;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (short)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("s", &objc_retval);
	return v;
}


/* signature: s16@4:8L12@16@20 */
static short 
meth_imp_602(id self, SEL sel, unsigned long arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	short objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("L", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("s", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_602(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	short objc_retval;
	unsigned long objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("L", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (short)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("s", &objc_retval);
	return v;
}


/* signature: s16@4:8r^{AEDesc=I^^{OpaqueAEDataStorageType}}12^{AEDesc=I^^{OpaqueAEDataStorageType}}16I20 */
static short 
meth_imp_603(id self, SEL sel, struct AEDesc  *arg_2, struct AEDesc  *arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	short objc_retval;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{AEDesc=I^^{OpaqueAEDataStorageType=}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{AEDesc=I^^{OpaqueAEDataStorageType=}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("s", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_603(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	short objc_retval;
	struct AEDesc  *objc_arg2;
	struct AEDesc  *objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{AEDesc=I^^{OpaqueAEDataStorageType=}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{AEDesc=I^^{OpaqueAEDataStorageType=}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (short)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("s", &objc_retval);
	return v;
}


/* signature: s4@4:8 */
static short 
meth_imp_604(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	short objc_retval;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("s", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_604(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	short objc_retval;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		objc_retval = (short)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("s", &objc_retval);
	return v;
}


/* signature: s8@4:8@12 */
static short 
meth_imp_605(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;
	const char* errstr;
	short objc_retval;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
	errstr = ObjC_PythonToObjC("s", retval, &objc_retval);
	Py_DECREF(retval);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_ValueError, "Cannot convert to ObjC");
		ObjCErr_ToObjC();
	}
	return objc_retval;
}
static PyObject* super_605(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	short objc_retval;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		objc_retval = (short)(long)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	v = ObjC_ObjCToPython("s", &objc_retval);
	return v;
}


/* signature: v104@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32{_NSRect={_NSPoint=ff}{_NSSize=ff}}48{_NSRect={_NSPoint=ff}{_NSSize=ff}}64{_NSRect={_NSPoint=ff}{_NSSize=ff}}80{_NSRect={_NSPoint=ff}{_NSSize=ff}}96 */
static void 
meth_imp_606(id self, SEL sel, struct _NSRect arg_2, struct _NSRect arg_3, struct _NSRect arg_4, struct _NSRect arg_5, struct _NSRect arg_6, struct _NSRect arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_606(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	struct _NSRect objc_arg3;
	struct _NSRect objc_arg4;
	struct _NSRect objc_arg5;
	struct _NSRect objc_arg6;
	struct _NSRect objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v10@4:8@12s16 */
static void 
meth_imp_607(id self, SEL sel, id arg_2, short arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_607(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	short objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v10@4:8^{OpaqueIconRef=}12s16 */
struct OpaqueIconRef;
static void 
meth_imp_608(id self, SEL sel, struct OpaqueIconRef  *arg_2, short arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{OpaqueIconRef=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("s", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_608(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaqueIconRef  *objc_arg2;
	short objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{OpaqueIconRef=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("s", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8#12^v16 */
static void 
meth_imp_609(id self, SEL sel, Class arg_2, void  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_609(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	Class objc_arg2;
	void  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8*12I16 */
static void 
meth_imp_610(id self, SEL sel, char* arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_610(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8:12@16 */
static void 
meth_imp_611(id self, SEL sel, SEL arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_611(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	SEL objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@12#16 */
static void 
meth_imp_612(id self, SEL sel, id arg_2, Class arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_612(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	Class objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@12:16 */
static void 
meth_imp_613(id self, SEL sel, id arg_2, SEL arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_613(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	SEL objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@12@16 */
static void 
meth_imp_614(id self, SEL sel, id arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_614(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@12I16 */
static void 
meth_imp_615(id self, SEL sel, id arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_615(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@12L16 */
static void 
meth_imp_616(id self, SEL sel, id arg_2, unsigned long arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("L", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_616(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	unsigned long objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("L", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@12^c16 */
static void 
meth_imp_617(id self, SEL sel, id arg_2, char  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_617(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	char  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@12^i16 */
static void 
meth_imp_618(id self, SEL sel, id arg_2, int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_618(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@12^v16 */
static void 
meth_imp_619(id self, SEL sel, id arg_2, void  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_619(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	void  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@12^{?=^SI^SI^SI}16 */
static void 
meth_imp_620(id self, SEL sel, id arg_2, struct pyobjcanonymous0  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_620(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct pyobjcanonymous0  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@12i16 */
static void 
meth_imp_621(id self, SEL sel, id arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_621(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@12l16 */
static void 
meth_imp_622(id self, SEL sel, id arg_2, long arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("l", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_622(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	long objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("l", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8@16 */
static void 
meth_imp_623(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_623(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8I12@16 */
static void 
meth_imp_624(id self, SEL sel, unsigned int arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_624(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8I12I16 */
static void 
meth_imp_625(id self, SEL sel, unsigned int arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_625(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8I12^v16 */
static void 
meth_imp_626(id self, SEL sel, unsigned int arg_2, void  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_626(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_arg2;
	void  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8Q12 */
static void 
meth_imp_627(id self, SEL sel, unsigned long long arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("Q", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_627(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned long long objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("Q", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8S12I16 */
static void 
meth_imp_628(id self, SEL sel, unsigned short arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_628(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned short objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^?12^v16 */
static void 
meth_imp_629(id self, SEL sel, void*  *arg_2, void  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^?", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_629(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void*  *objc_arg2;
	void  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^?", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^@12^@16 */
static void 
meth_imp_630(id self, SEL sel, id  *arg_2, id  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_630(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id  *objc_arg2;
	id  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^@12^i16 */
static void 
meth_imp_631(id self, SEL sel, id  *arg_2, int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_631(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id  *objc_arg2;
	int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^@12^{_NSRange=II}16 */
static void 
meth_imp_632(id self, SEL sel, id  *arg_2, struct _NSRange  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_632(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id  *objc_arg2;
	struct _NSRange  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^@12^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
static void 
meth_imp_633(id self, SEL sel, id  *arg_2, struct _NSRect  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_633(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id  *objc_arg2;
	struct _NSRect  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^I12I16 */
static void 
meth_imp_634(id self, SEL sel, unsigned int  *arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_634(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int  *objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^I12^I16 */
static void 
meth_imp_635(id self, SEL sel, unsigned int  *arg_2, unsigned int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_635(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int  *objc_arg2;
	unsigned int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^^S12^i16 */
static void 
meth_imp_636(id self, SEL sel, unsigned short  * *arg_2, int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^^S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_636(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned short  * *objc_arg2;
	int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^^S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^^{OpaqueIconRef}12^s16 */
struct OpaqueIconRef;
static void 
meth_imp_637(id self, SEL sel, struct OpaqueIconRef  * *arg_2, short  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^^{OpaqueIconRef=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^s", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_637(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaqueIconRef  * *objc_arg2;
	short  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^^{OpaqueIconRef=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^s", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^f12^f16 */
static void 
meth_imp_638(id self, SEL sel, float  *arg_2, float  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_638(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float  *objc_arg2;
	float  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^i12I16 */
static void 
meth_imp_639(id self, SEL sel, int  *arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_639(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^i12^f16 */
static void 
meth_imp_640(id self, SEL sel, int  *arg_2, float  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_640(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_arg2;
	float  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^i12^i16 */
static void 
meth_imp_641(id self, SEL sel, int  *arg_2, int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_641(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_arg2;
	int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^l12i16 */
static void 
meth_imp_642(id self, SEL sel, long  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^l", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_642(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	long  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^l", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^v12I16 */
static void 
meth_imp_643(id self, SEL sel, void  *arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_643(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^v12i16 */
static void 
meth_imp_644(id self, SEL sel, void  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_644(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^{_NSPoint=ff}12i16 */
static void 
meth_imp_645(id self, SEL sel, struct _NSPoint  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_645(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12i16 */
static void 
meth_imp_646(id self, SEL sel, struct _NSRect  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_646(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}12i16 */
struct _RowEntry;
static void 
meth_imp_647(id self, SEL sel, struct _RowEntry  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_RowEntry=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_647(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _RowEntry  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_RowEntry=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8^{__CFReadStream=}12@16 */
struct __CFReadStream;
static void 
meth_imp_648(id self, SEL sel, struct __CFReadStream  *arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{__CFReadStream=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_648(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFReadStream  *objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{__CFReadStream=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8c12@16 */
static void 
meth_imp_649(id self, SEL sel, char arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_649(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8c12I16 */
static void 
meth_imp_650(id self, SEL sel, char arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_650(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8i12@16 */
static void 
meth_imp_651(id self, SEL sel, int arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_651(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8i12I16 */
static void 
meth_imp_652(id self, SEL sel, int arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_652(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8i12i16 */
static void 
meth_imp_653(id self, SEL sel, int arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_653(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8r*12^v16 */
static void 
meth_imp_654(id self, SEL sel, char* arg_2, void  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_654(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_arg2;
	void  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8r*12i16 */
static void 
meth_imp_655(id self, SEL sel, char* arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_655(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8r*12r^v16 */
static void 
meth_imp_656(id self, SEL sel, char* arg_2, void  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_656(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_arg2;
	void  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8r*16 */
static void 
meth_imp_657(id self, SEL sel, char* arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_657(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8r^S12i16 */
static void 
meth_imp_658(id self, SEL sel, unsigned short  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_658(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned short  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8r^^i12^i16 */
static void 
meth_imp_659(id self, SEL sel, int  * *arg_2, int  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_659(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  * *objc_arg2;
	int  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8r^i12i16 */
static void 
meth_imp_660(id self, SEL sel, int  *arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_660(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8r^v12I16 */
static void 
meth_imp_661(id self, SEL sel, void  *arg_2, unsigned int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_661(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	unsigned int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8r^{_NSPoint=ff}12@16 */
static void 
meth_imp_662(id self, SEL sel, struct _NSPoint  *arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_662(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint  *objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8{_NSPoint=ff}12 */
static void 
meth_imp_663(id self, SEL sel, struct _NSPoint arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_663(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8{_NSRange=II}12 */
static void 
meth_imp_664(id self, SEL sel, struct _NSRange arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_664(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v12@4:8{_NSSize=ff}12 */
static void 
meth_imp_665(id self, SEL sel, struct _NSSize arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_665(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSSize objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v13@4:8:12@16c20 */
static void 
meth_imp_666(id self, SEL sel, SEL arg_2, id arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_666(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	SEL objc_arg2;
	id objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v13@4:8@12@16c20 */
static void 
meth_imp_667(id self, SEL sel, id arg_2, id arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_667(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v13@4:8@12^i16c20 */
static void 
meth_imp_668(id self, SEL sel, id arg_2, int  *arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_668(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int  *objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v13@4:8@12c16c20 */
static void 
meth_imp_669(id self, SEL sel, id arg_2, char arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_669(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	char objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v13@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@16c20 */
static void 
meth_imp_670(id self, SEL sel, struct _NSRect  *arg_2, id arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_670(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect  *objc_arg2;
	id objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v13@4:8i12c16c20 */
static void 
meth_imp_671(id self, SEL sel, int arg_2, char arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_671(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	char objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v13@4:8i12i16c20 */
static void 
meth_imp_672(id self, SEL sel, int arg_2, int arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_672(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	int objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v13@4:8{_NSRange=II}12c20 */
static void 
meth_imp_673(id self, SEL sel, struct _NSRange arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_673(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8:12@16@20 */
static void 
meth_imp_674(id self, SEL sel, SEL arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_674(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	SEL objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8:12i16i20 */
static void 
meth_imp_675(id self, SEL sel, SEL arg_2, int arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_675(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	SEL objc_arg2;
	int objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12:16#20 */
static void 
meth_imp_676(id self, SEL sel, id arg_2, SEL arg_3, Class arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_676(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	SEL objc_arg3;
	Class objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12:16@20 */
static void 
meth_imp_677(id self, SEL sel, id arg_2, SEL arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_677(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	SEL objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12:16I20 */
static void 
meth_imp_678(id self, SEL sel, id arg_2, SEL arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_678(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	SEL objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12:16^v20 */
static void 
meth_imp_679(id self, SEL sel, id arg_2, SEL arg_3, void  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_679(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	SEL objc_arg3;
	void  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12@16*20 */
static void 
meth_imp_680(id self, SEL sel, id arg_2, id arg_3, char* arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_680(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	char* objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12@16@20 */
static void 
meth_imp_681(id self, SEL sel, id arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_681(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12@16I20 */
static void 
meth_imp_682(id self, SEL sel, id arg_2, id arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_682(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12@16L20 */
static void 
meth_imp_683(id self, SEL sel, id arg_2, id arg_3, unsigned long arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("L", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_683(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	unsigned long objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("L", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12@16i20 */
static void 
meth_imp_684(id self, SEL sel, id arg_2, id arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_684(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12@20 */
static void 
meth_imp_685(id self, SEL sel, id arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_685(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12I16@20 */
static void 
meth_imp_686(id self, SEL sel, id arg_2, unsigned int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_686(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	unsigned int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12^@16^@20 */
static void 
meth_imp_687(id self, SEL sel, id arg_2, id  *arg_3, id  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_687(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id  *objc_arg3;
	id  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12c16^v20 */
static void 
meth_imp_688(id self, SEL sel, id arg_2, char arg_3, void  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_688(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	char objc_arg3;
	void  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12i16@20 */
static void 
meth_imp_689(id self, SEL sel, id arg_2, int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_689(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12i16I20 */
static void 
meth_imp_690(id self, SEL sel, id arg_2, int arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_690(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12i16^v20 */
static void 
meth_imp_691(id self, SEL sel, id arg_2, int arg_3, void  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_691(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	void  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12i16i20 */
static void 
meth_imp_692(id self, SEL sel, id arg_2, int arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_692(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12{_NSPoint=ff}16 */
static void 
meth_imp_693(id self, SEL sel, id arg_2, struct _NSPoint arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_693(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSPoint objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12{_NSRange=II}16 */
static void 
meth_imp_694(id self, SEL sel, id arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_694(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8@12{_NSSize=ff}16 */
static void 
meth_imp_695(id self, SEL sel, id arg_2, struct _NSSize arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_695(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSSize objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8I12@16@20 */
static void 
meth_imp_696(id self, SEL sel, unsigned int arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_696(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8I12I16I20 */
static void 
meth_imp_697(id self, SEL sel, unsigned int arg_2, unsigned int arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_697(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_arg2;
	unsigned int objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8I12^v16L20 */
static void 
meth_imp_698(id self, SEL sel, unsigned int arg_2, void  *arg_3, unsigned long arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("L", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_698(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_arg2;
	void  *objc_arg3;
	unsigned long objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("L", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^@12{_NSRange=II}16 */
static void 
meth_imp_699(id self, SEL sel, id  *arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_699(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id  *objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^I12i16@20 */
static void 
meth_imp_700(id self, SEL sel, unsigned int  *arg_2, int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_700(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int  *objc_arg2;
	int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^S12^i16^{?=^SI^SI^SI}20 */
static void 
meth_imp_701(id self, SEL sel, unsigned short  *arg_2, int  *arg_3, struct pyobjcanonymous0  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_701(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned short  *objc_arg2;
	int  *objc_arg3;
	struct pyobjcanonymous0  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^S12{_NSRange=II}16 */
static void 
meth_imp_702(id self, SEL sel, unsigned short  *arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_702(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned short  *objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^^{OpaqueIconRef}12^s16@20 */
struct OpaqueIconRef;
static void 
meth_imp_703(id self, SEL sel, struct OpaqueIconRef  * *arg_2, short  *arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^^{OpaqueIconRef=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^s", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_703(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaqueIconRef  * *objc_arg2;
	short  *objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^^{OpaqueIconRef=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^s", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^f12^i16^f20 */
static void 
meth_imp_704(id self, SEL sel, float  *arg_2, int  *arg_3, float  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_704(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float  *objc_arg2;
	int  *objc_arg3;
	float  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^i12I16I20 */
static void 
meth_imp_705(id self, SEL sel, int  *arg_2, unsigned int arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_705(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_arg2;
	unsigned int objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^i12I16^I20 */
static void 
meth_imp_706(id self, SEL sel, int  *arg_2, unsigned int arg_3, unsigned int  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_706(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_arg2;
	unsigned int objc_arg3;
	unsigned int  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^l12i16i20 */
static void 
meth_imp_707(id self, SEL sel, long  *arg_2, int arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^l", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_707(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	long  *objc_arg2;
	int objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^l", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^v12I16I20 */
static void 
meth_imp_708(id self, SEL sel, void  *arg_2, unsigned int arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_708(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	unsigned int objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^v12I16^I20 */
static void 
meth_imp_709(id self, SEL sel, void  *arg_2, unsigned int arg_3, unsigned int  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_709(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	unsigned int objc_arg3;
	unsigned int  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^v12{_NSRange=II}16 */
static void 
meth_imp_710(id self, SEL sel, void  *arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_710(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^{_NSMapTable=}12r*16@20 */
struct _NSMapTable;
static void 
meth_imp_711(id self, SEL sel, struct _NSMapTable  *arg_2, char* arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSMapTable=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_711(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSMapTable  *objc_arg2;
	char* objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSMapTable=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^{__CFData=}12^{__CFData=}16^{__CFSocket=}20 */
struct __CFData;
struct __CFData;
struct __CFSocket;
static void 
meth_imp_712(id self, SEL sel, struct __CFData  *arg_2, struct __CFData  *arg_3, struct __CFSocket  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{__CFData=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{__CFData=}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{__CFSocket=}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_712(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFData  *objc_arg2;
	struct __CFData  *objc_arg3;
	struct __CFSocket  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{__CFData=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{__CFData=}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{__CFSocket=}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8^{__CFString=}12I16I20 */
struct __CFString;
static void 
meth_imp_713(id self, SEL sel, struct __CFString  *arg_2, unsigned int arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{__CFString=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_713(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFString  *objc_arg2;
	unsigned int objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{__CFString=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8c12I16I20 */
static void 
meth_imp_714(id self, SEL sel, char arg_2, unsigned int arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_714(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	unsigned int objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8c12i16i20 */
static void 
meth_imp_715(id self, SEL sel, char arg_2, int arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_715(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	int objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8c12{_NSPoint=ff}16 */
static void 
meth_imp_716(id self, SEL sel, char arg_2, struct _NSPoint arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_716(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	struct _NSPoint objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8i12Q16 */
static void 
meth_imp_717(id self, SEL sel, int arg_2, unsigned long long arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("Q", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_717(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	unsigned long long objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("Q", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8i12i16@20 */
static void 
meth_imp_718(id self, SEL sel, int arg_2, int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_718(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8i12i16I20 */
static void 
meth_imp_719(id self, SEL sel, int arg_2, int arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_719(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	int objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8i12i16i20 */
static void 
meth_imp_720(id self, SEL sel, int arg_2, int arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_720(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	int objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8i12{_NSRange=II}16 */
static void 
meth_imp_721(id self, SEL sel, int arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_721(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8q12@20 */
static void 
meth_imp_722(id self, SEL sel, long long arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("q", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_722(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	long long objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("q", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8r*12I16^v20 */
static void 
meth_imp_723(id self, SEL sel, char* arg_2, unsigned int arg_3, void  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_723(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_arg2;
	unsigned int objc_arg3;
	void  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8r*12I16r^v20 */
static void 
meth_imp_724(id self, SEL sel, char* arg_2, unsigned int arg_3, void  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_724(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_arg2;
	unsigned int objc_arg3;
	void  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8r*12{_NSPoint=ff}16 */
static void 
meth_imp_725(id self, SEL sel, char* arg_2, struct _NSPoint arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_725(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_arg2;
	struct _NSPoint objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8{_NSPoint=ff}12@20 */
static void 
meth_imp_726(id self, SEL sel, struct _NSPoint arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_726(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8{_NSPoint=ff}12i20 */
static void 
meth_imp_727(id self, SEL sel, struct _NSPoint arg_2, int arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_727(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	int objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8{_NSRange=II}12@20 */
static void 
meth_imp_728(id self, SEL sel, struct _NSRange arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_728(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v16@4:8{_NSRange=II}12r^v20 */
static void 
meth_imp_729(id self, SEL sel, struct _NSRange arg_2, void  *arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_729(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	void  *objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v17@4:8@12@16@20c24 */
static void 
meth_imp_730(id self, SEL sel, id arg_2, id arg_3, id arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_730(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v17@4:8@12c16c20c24 */
static void 
meth_imp_731(id self, SEL sel, id arg_2, char arg_3, char arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_731(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	char objc_arg3;
	char objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v17@4:8@12{_NSRange=II}16c24 */
static void 
meth_imp_732(id self, SEL sel, id arg_2, struct _NSRange arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_732(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSRange objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v17@4:8^v12I16c20c24 */
static void 
meth_imp_733(id self, SEL sel, void  *arg_2, unsigned int arg_3, char arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_733(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	unsigned int objc_arg3;
	char objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v17@4:8^v12{_NSRange=II}16c24 */
static void 
meth_imp_734(id self, SEL sel, void  *arg_2, struct _NSRange arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_734(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	struct _NSRange objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v17@4:8i12c16c20c24 */
static void 
meth_imp_735(id self, SEL sel, int arg_2, char arg_3, char arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_735(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	char objc_arg3;
	char objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v17@4:8i12i16@20c24 */
static void 
meth_imp_736(id self, SEL sel, int arg_2, int arg_3, id arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_736(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	int objc_arg3;
	id objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v17@4:8i12i16i20c24 */
static void 
meth_imp_737(id self, SEL sel, int arg_2, int arg_3, int arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_737(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	int objc_arg3;
	int objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v17@4:8{_NSRange=II}12^v20c24 */
static void 
meth_imp_738(id self, SEL sel, struct _NSRange arg_2, void  *arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_738(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	void  *objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v17@4:8{_NSRange=II}12i20c24 */
static void 
meth_imp_739(id self, SEL sel, struct _NSRange arg_2, int arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_739(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	int objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12:16#20#24 */
static void 
meth_imp_740(id self, SEL sel, id arg_2, SEL arg_3, Class arg_4, Class arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_740(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	SEL objc_arg3;
	Class objc_arg4;
	Class objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12:16@20@24 */
static void 
meth_imp_741(id self, SEL sel, id arg_2, SEL arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_741(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	SEL objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12:16I20I24 */
static void 
meth_imp_742(id self, SEL sel, id arg_2, SEL arg_3, unsigned int arg_4, unsigned int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_742(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	SEL objc_arg3;
	unsigned int objc_arg4;
	unsigned int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12@16:20^v24 */
static void 
meth_imp_743(id self, SEL sel, id arg_2, id arg_3, SEL arg_4, void  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_743(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	SEL objc_arg4;
	void  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12@16@20@24 */
static void 
meth_imp_744(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_744(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12@16@20I24 */
static void 
meth_imp_745(id self, SEL sel, id arg_2, id arg_3, id arg_4, unsigned int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_745(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	unsigned int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12@16@20i24 */
static void 
meth_imp_746(id self, SEL sel, id arg_2, id arg_3, id arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_746(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12@16I20@24 */
static void 
meth_imp_747(id self, SEL sel, id arg_2, id arg_3, unsigned int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_747(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12@16i20@24 */
static void 
meth_imp_748(id self, SEL sel, id arg_2, id arg_3, int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_748(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12@16i20i24 */
static void 
meth_imp_749(id self, SEL sel, id arg_2, id arg_3, int arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_749(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12@16l20@24 */
static void 
meth_imp_750(id self, SEL sel, id arg_2, id arg_3, long arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("l", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_750(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	long objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("l", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12@16{_NSRange=II}20 */
static void 
meth_imp_751(id self, SEL sel, id arg_2, id arg_3, struct _NSRange arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_751(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	struct _NSRange objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12I16@20*24 */
static void 
meth_imp_752(id self, SEL sel, id arg_2, unsigned int arg_3, id arg_4, char* arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_752(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	unsigned int objc_arg3;
	id objc_arg4;
	char* objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12I16@24 */
static void 
meth_imp_753(id self, SEL sel, id arg_2, unsigned int arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_753(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	unsigned int objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12I16I20^I24 */
static void 
meth_imp_754(id self, SEL sel, id arg_2, unsigned int arg_3, unsigned int arg_4, unsigned int  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_754(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	unsigned int objc_arg3;
	unsigned int objc_arg4;
	unsigned int  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12^{__CFPasteboard=}16i20^v24 */
struct __CFPasteboard;
static void 
meth_imp_755(id self, SEL sel, id arg_2, struct __CFPasteboard  *arg_3, int arg_4, void  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{__CFPasteboard=}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_755(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct __CFPasteboard  *objc_arg3;
	int objc_arg4;
	void  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{__CFPasteboard=}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12c16i20i24 */
static void 
meth_imp_756(id self, SEL sel, id arg_2, char arg_3, int arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_756(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	char objc_arg3;
	int objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12i16I20@24 */
static void 
meth_imp_757(id self, SEL sel, id arg_2, int arg_3, unsigned int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_757(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	unsigned int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12{_NSPoint=ff}16I24 */
static void 
meth_imp_758(id self, SEL sel, id arg_2, struct _NSPoint arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_758(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSPoint objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8@12{_NSRange=II}16@24 */
static void 
meth_imp_759(id self, SEL sel, id arg_2, struct _NSRange arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_759(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSRange objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8I12{_NSRange=II}16i24 */
static void 
meth_imp_760(id self, SEL sel, unsigned int arg_2, struct _NSRange arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_760(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_arg2;
	struct _NSRange objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8^?12^v16{_NSRange=II}20 */
static void 
meth_imp_761(id self, SEL sel, void*  *arg_2, void  *arg_3, struct _NSRange arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^?", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_761(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void*  *objc_arg2;
	void  *objc_arg3;
	struct _NSRange objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^?", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8^f12^f16^f20^f24 */
static void 
meth_imp_762(id self, SEL sel, float  *arg_2, float  *arg_3, float  *arg_4, float  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_762(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float  *objc_arg2;
	float  *objc_arg3;
	float  *objc_arg4;
	float  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8^i12^i16{_NSPoint=ff}20 */
static void 
meth_imp_763(id self, SEL sel, int  *arg_2, int  *arg_3, struct _NSPoint arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_763(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_arg2;
	int  *objc_arg3;
	struct _NSPoint objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8^v12l16l20l24 */
static void 
meth_imp_764(id self, SEL sel, void  *arg_2, long arg_3, long arg_4, long arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("l", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("l", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("l", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_764(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	long objc_arg3;
	long objc_arg4;
	long objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("l", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("l", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("l", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8^v12r*16^I20@24 */
static void 
meth_imp_765(id self, SEL sel, void  *arg_2, char* arg_3, unsigned int  *arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_765(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	char* objc_arg3;
	unsigned int  *objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8c12@16@20@24 */
static void 
meth_imp_766(id self, SEL sel, char arg_2, id arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_766(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8i12@16:20^v24 */
static void 
meth_imp_767(id self, SEL sel, int arg_2, id arg_3, SEL arg_4, void  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_767(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	id objc_arg3;
	SEL objc_arg4;
	void  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSPoint=ff}12{_NSPoint=ff}20 */
static void 
meth_imp_768(id self, SEL sel, struct _NSPoint arg_2, struct _NSPoint arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_768(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	struct _NSPoint objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSPoint=ff}12{_NSRange=II}20 */
static void 
meth_imp_769(id self, SEL sel, struct _NSPoint arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_769(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSRange=II}12@20I24 */
static void 
meth_imp_770(id self, SEL sel, struct _NSRange arg_2, id arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_770(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSRange=II}12^@20I24 */
static void 
meth_imp_771(id self, SEL sel, struct _NSRange arg_2, id  *arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_771(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	id  *objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSRange=II}12c20^{_NSRange=II}24 */
static void 
meth_imp_772(id self, SEL sel, struct _NSRange arg_2, char arg_3, struct _NSRange  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_772(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	char objc_arg3;
	struct _NSRange  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSRange=II}12i20^{_NSRange=II}24 */
static void 
meth_imp_773(id self, SEL sel, struct _NSRange arg_2, int arg_3, struct _NSRange  *arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_773(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	int objc_arg3;
	struct _NSRange  *objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSRange=II}12r*20I24 */
static void 
meth_imp_774(id self, SEL sel, struct _NSRange arg_2, char* arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_774(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	char* objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSRange=II}12r^S20I24 */
static void 
meth_imp_775(id self, SEL sel, struct _NSRange arg_2, unsigned short  *arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^S", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_775(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	unsigned short  *objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^S", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSRange=II}12{_NSRange=II}20 */
static void 
meth_imp_776(id self, SEL sel, struct _NSRange arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_776(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12 */
static void 
meth_imp_777(id self, SEL sel, struct _NSRect arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_777(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSSize=ff}12{_NSRange=II}20 */
static void 
meth_imp_778(id self, SEL sel, struct _NSSize arg_2, struct _NSRange arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_778(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSSize objc_arg2;
	struct _NSRange objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v20@4:8{_NSSize=ff}12{_NSSize=ff}20 */
static void 
meth_imp_779(id self, SEL sel, struct _NSSize arg_2, struct _NSSize arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_779(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSSize objc_arg2;
	struct _NSSize objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v21@4:8@12@16@20@24c28 */
static void 
meth_imp_780(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_780(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v21@4:8@12i16c20c24c28 */
static void 
meth_imp_781(id self, SEL sel, id arg_2, int arg_3, char arg_4, char arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_781(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	char objc_arg4;
	char objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v21@4:8@12i16i20i24c28 */
static void 
meth_imp_782(id self, SEL sel, id arg_2, int arg_3, int arg_4, int arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_782(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	int objc_arg4;
	int objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v21@4:8i12i16c20c24c28 */
static void 
meth_imp_783(id self, SEL sel, int arg_2, int arg_3, char arg_4, char arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_783(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	int objc_arg3;
	char objc_arg4;
	char objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v21@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28 */
static void 
meth_imp_784(id self, SEL sel, struct _NSRect arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_784(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8*12I16{_NSRange=II}20^{_NSRange=II}28 */
static void 
meth_imp_785(id self, SEL sel, char* arg_2, unsigned int arg_3, struct _NSRange arg_4, struct _NSRange  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_785(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_arg2;
	unsigned int objc_arg3;
	struct _NSRange objc_arg4;
	struct _NSRange  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8:12@16@20I24@28 */
static void 
meth_imp_786(id self, SEL sel, SEL arg_2, id arg_3, id arg_4, unsigned int arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_786(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	SEL objc_arg2;
	id objc_arg3;
	id objc_arg4;
	unsigned int objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8@12:16@20@24I28 */
static void 
meth_imp_787(id self, SEL sel, id arg_2, SEL arg_3, id arg_4, id arg_5, unsigned int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_787(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	SEL objc_arg3;
	id objc_arg4;
	id objc_arg5;
	unsigned int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8@12:16@20@24i28 */
static void 
meth_imp_788(id self, SEL sel, id arg_2, SEL arg_3, id arg_4, id arg_5, int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_788(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	SEL objc_arg3;
	id objc_arg4;
	id objc_arg5;
	int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8@12@16@20:24^v28 */
static void 
meth_imp_789(id self, SEL sel, id arg_2, id arg_3, id arg_4, SEL arg_5, void  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_789(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	SEL objc_arg5;
	void  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8@12@16@20I24@28 */
static void 
meth_imp_790(id self, SEL sel, id arg_2, id arg_3, id arg_4, unsigned int arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_790(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	unsigned int objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8@12@16i20@28 */
static void 
meth_imp_791(id self, SEL sel, id arg_2, id arg_3, int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_791(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8@12c16@20:24^v28 */
static void 
meth_imp_792(id self, SEL sel, id arg_2, char arg_3, id arg_4, SEL arg_5, void  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_792(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	char objc_arg3;
	id objc_arg4;
	SEL objc_arg5;
	void  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8@12i16@20:24^v28 */
static void 
meth_imp_793(id self, SEL sel, id arg_2, int arg_3, id arg_4, SEL arg_5, void  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_793(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	id objc_arg4;
	SEL objc_arg5;
	void  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8@12{_NSPoint=ff}16{_NSPoint=ff}24 */
static void 
meth_imp_794(id self, SEL sel, id arg_2, struct _NSPoint arg_3, struct _NSPoint arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_794(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSPoint objc_arg3;
	struct _NSPoint objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8@12{_NSRange=II}16{_NSRange=II}24 */
static void 
meth_imp_795(id self, SEL sel, id arg_2, struct _NSRange arg_3, struct _NSRange arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_795(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSRange objc_arg3;
	struct _NSRange objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
static void 
meth_imp_796(id self, SEL sel, id arg_2, struct _NSRect arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_796(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSRect objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8I12{_NSPoint=ff}16I24@28 */
static void 
meth_imp_797(id self, SEL sel, unsigned int arg_2, struct _NSPoint arg_3, unsigned int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_797(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_arg2;
	struct _NSPoint objc_arg3;
	unsigned int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8^I12^I16^I20{_NSRange=II}24 */
static void 
meth_imp_798(id self, SEL sel, unsigned int  *arg_2, unsigned int  *arg_3, unsigned int  *arg_4, struct _NSRange arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_798(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int  *objc_arg2;
	unsigned int  *objc_arg3;
	unsigned int  *objc_arg4;
	struct _NSRange objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8^f12^f16^f20^f24^f28 */
static void 
meth_imp_799(id self, SEL sel, float  *arg_2, float  *arg_3, float  *arg_4, float  *arg_5, float  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_799(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float  *objc_arg2;
	float  *objc_arg3;
	float  *objc_arg4;
	float  *objc_arg5;
	float  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8^v12^@16^@20^I24^@28 */
static void 
meth_imp_800(id self, SEL sel, void  *arg_2, id  *arg_3, id  *arg_4, unsigned int  *arg_5, id  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_800(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	id  *objc_arg3;
	id  *objc_arg4;
	unsigned int  *objc_arg5;
	id  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8^{_NSGlyphGenContext=iiiiiiiiiii@[32i][32i][32i][64i]{_NSRange=II}{_NSRange=II}ii^{_NSGlyphInsertBuffer}}12@16@20^{_NSRAStringBuffer=@IIIIII[100S]}24@28 */
struct _NSGlyphInsertBuffer;struct _NSGlyphGenContext {
	int field_0;
	int field_1;
	int field_2;
	int field_3;
	int field_4;
	int field_5;
	int field_6;
	int field_7;
	int field_8;
	int field_9;
	int field_10;
	id field_11;
	int field_12[32];
	int field_13[32];
	int field_14[32];
	int field_15[64];
	struct _NSRange field_16;
	struct _NSRange field_17;
	int field_18;
	int field_19;
	struct _NSGlyphInsertBuffer  *field_20;
};

struct _NSRAStringBuffer {
	id field_0;
	unsigned int field_1;
	unsigned int field_2;
	unsigned int field_3;
	unsigned int field_4;
	unsigned int field_5;
	unsigned int field_6;
	unsigned short field_7[100];
};

static void 
meth_imp_801(id self, SEL sel, struct _NSGlyphGenContext  *arg_2, id arg_3, id arg_4, struct _NSRAStringBuffer  *arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSGlyphGenContext=iiiiiiiiiii@[32i][32i][32i][64i]{_NSRange=II}{_NSRange=II}ii^{_NSGlyphInsertBuffer=}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRAStringBuffer=@IIIIII[100S]}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_801(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSGlyphGenContext  *objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct _NSRAStringBuffer  *objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSGlyphGenContext=iiiiiiiiiii@[32i][32i][32i][64i]{_NSRange=II}{_NSRange=II}ii^{_NSGlyphInsertBuffer=}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSRAStringBuffer=@IIIIII[100S]}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
static void 
meth_imp_802(id self, SEL sel, struct _NSRect  *arg_2, struct _NSRect arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_802(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect  *objc_arg2;
	struct _NSRect objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8c12I16r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}20r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}24^{_NSRect={_NSPoint=ff}{_NSSize=ff}}28 */
static void 
meth_imp_803(id self, SEL sel, char arg_2, unsigned int arg_3, struct _NSRect  *arg_4, struct _NSRect  *arg_5, struct _NSRect  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_803(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	unsigned int objc_arg3;
	struct _NSRect  *objc_arg4;
	struct _NSRect  *objc_arg5;
	struct _NSRect  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8c12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
static void 
meth_imp_804(id self, SEL sel, char arg_2, struct _NSRect arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_804(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	struct _NSRect objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8i12@16:20i24i28 */
static void 
meth_imp_805(id self, SEL sel, int arg_2, id arg_3, SEL arg_4, int arg_5, int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_805(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	id objc_arg3;
	SEL objc_arg4;
	int objc_arg5;
	int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8i12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16 */
static void 
meth_imp_806(id self, SEL sel, int arg_2, struct _NSRect arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_806(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	struct _NSRect objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8{_NSPoint=ff}12{_NSPoint=ff}20@28 */
static void 
meth_imp_807(id self, SEL sel, struct _NSPoint arg_2, struct _NSPoint arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_807(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	struct _NSPoint objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8{_NSRange=II}12@20{_NSRange=II}24 */
static void 
meth_imp_808(id self, SEL sel, struct _NSRange arg_2, id arg_3, struct _NSRange arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_808(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	id objc_arg3;
	struct _NSRange objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28 */
static void 
meth_imp_809(id self, SEL sel, struct _NSRect arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_809(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v24@4:8{_NSSize=ff}12^{_NSSize=ff}20^{_NSRect={_NSPoint=ff}{_NSSize=ff}}24^{_NSRect={_NSPoint=ff}{_NSSize=ff}}28 */
static void 
meth_imp_810(id self, SEL sel, struct _NSSize arg_2, struct _NSSize  *arg_3, struct _NSRect  *arg_4, struct _NSRect  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSSize=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_810(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSSize objc_arg2;
	struct _NSSize  *objc_arg3;
	struct _NSRect  *objc_arg4;
	struct _NSRect  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSSize=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v25@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16c32 */
static void 
meth_imp_811(id self, SEL sel, id arg_2, struct _NSRect arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_811(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSRect objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v25@4:8i12i16c20c24c28c32 */
static void 
meth_imp_812(id self, SEL sel, int arg_2, int arg_3, char arg_4, char arg_5, char arg_6, char arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_812(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	int objc_arg3;
	char objc_arg4;
	char objc_arg5;
	char objc_arg6;
	char objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v25@4:8{_NSPoint=ff}12{_NSPoint=ff}20@28c32 */
static void 
meth_imp_813(id self, SEL sel, struct _NSPoint arg_2, struct _NSPoint arg_3, id arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_813(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	struct _NSPoint objc_arg3;
	id objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v25@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28c32 */
static void 
meth_imp_814(id self, SEL sel, struct _NSRect arg_2, id arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_814(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	id objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v25@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28c32 */
static void 
meth_imp_815(id self, SEL sel, struct _NSRect arg_2, char arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_815(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	char objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8:12@16@20i24@32 */
static void 
meth_imp_816(id self, SEL sel, SEL arg_2, id arg_3, id arg_4, int arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_816(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	SEL objc_arg2;
	id objc_arg3;
	id objc_arg4;
	int objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8@12@16@20@24:28^v32 */
static void 
meth_imp_817(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, SEL arg_6, void  *arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_817(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	SEL objc_arg6;
	void  *objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8@12@16i20@24:28^v32 */
static void 
meth_imp_818(id self, SEL sel, id arg_2, id arg_3, int arg_4, id arg_5, SEL arg_6, void  *arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_818(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	int objc_arg4;
	id objc_arg5;
	SEL objc_arg6;
	void  *objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8@12@16{_NSRect={_NSPoint=ff}{_NSSize=ff}}20 */
static void 
meth_imp_819(id self, SEL sel, id arg_2, id arg_3, struct _NSRect arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_819(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	struct _NSRect objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8@12i16{_NSRect={_NSPoint=ff}{_NSSize=ff}}20 */
static void 
meth_imp_820(id self, SEL sel, id arg_2, int arg_3, struct _NSRect arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_820(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	struct _NSRect objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32 */
static void 
meth_imp_821(id self, SEL sel, id arg_2, struct _NSRect arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_821(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8@12{_NSSize=ff}16i24^i28^i32 */
static void 
meth_imp_822(id self, SEL sel, id arg_2, struct _NSSize arg_3, int arg_4, int  *arg_5, int  *arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_822(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSSize objc_arg3;
	int objc_arg4;
	int  *objc_arg5;
	int  *objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8I12{_NSRange=II}16i24{_NSRange=II}28 */
static void 
meth_imp_823(id self, SEL sel, unsigned int arg_2, struct _NSRange arg_3, int arg_4, struct _NSRange arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_823(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_arg2;
	struct _NSRange objc_arg3;
	int objc_arg4;
	struct _NSRange objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8^{_PartStruct=if}12^I16{_NSRect={_NSPoint=ff}{_NSSize=ff}}20 */
struct _PartStruct {
	int field_0;
	float field_1;
};

static void 
meth_imp_824(id self, SEL sel, struct _PartStruct  *arg_2, unsigned int  *arg_3, struct _NSRect arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_PartStruct=if}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_824(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _PartStruct  *objc_arg2;
	unsigned int  *objc_arg3;
	struct _NSRect objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_PartStruct=if}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8c12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32 */
static void 
meth_imp_825(id self, SEL sel, char arg_2, struct _NSRect arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_825(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8i12^{_NSGlyphGenContext=iiiiiiiiiii@[32i][32i][32i][64i]{_NSRange=II}{_NSRange=II}ii^{_NSGlyphInsertBuffer}}16@20@24^{_NSRAStringBuffer=@IIIIII[100S]}28@32 */
static void 
meth_imp_826(id self, SEL sel, int arg_2, struct _NSGlyphGenContext  *arg_3, id arg_4, id arg_5, struct _NSRAStringBuffer  *arg_6, id arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^{_NSGlyphGenContext=iiiiiiiiiii@[32i][32i][32i][64i]{_NSRange=II}{_NSRange=II}ii^{_NSGlyphInsertBuffer=}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRAStringBuffer=@IIIIII[100S]}", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_826(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	struct _NSGlyphGenContext  *objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct _NSRAStringBuffer  *objc_arg6;
	id objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^{_NSGlyphGenContext=iiiiiiiiiii@[32i][32i][32i][64i]{_NSRange=II}{_NSRange=II}ii^{_NSGlyphInsertBuffer=}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^{_NSRAStringBuffer=@IIIIII[100S]}", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8{_NSAffineTransformStruct=ffffff}12 */
struct _NSAffineTransformStruct {
	float field_0;
	float field_1;
	float field_2;
	float field_3;
	float field_4;
	float field_5;
};

static void 
meth_imp_827(id self, SEL sel, struct _NSAffineTransformStruct arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSAffineTransformStruct=ffffff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_827(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSAffineTransformStruct objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSAffineTransformStruct=ffffff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8{_NSPoint=ff}12{_NSPoint=ff}20{_NSPoint=ff}28 */
static void 
meth_imp_828(id self, SEL sel, struct _NSPoint arg_2, struct _NSPoint arg_3, struct _NSPoint arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_828(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	struct _NSPoint objc_arg3;
	struct _NSPoint objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8{_NSRange=II}12{_NSRange=II}20i28^{_NSRange=II}32 */
static void 
meth_imp_829(id self, SEL sel, struct _NSRange arg_2, struct _NSRange arg_3, int arg_4, struct _NSRange  *arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_829(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRange objc_arg2;
	struct _NSRange objc_arg3;
	int objc_arg4;
	struct _NSRange  *objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32 */
static void 
meth_imp_830(id self, SEL sel, struct _NSRect arg_2, id arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_830(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	id objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28I32 */
static void 
meth_imp_831(id self, SEL sel, struct _NSRect arg_2, id arg_3, unsigned int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_831(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28@32 */
static void 
meth_imp_832(id self, SEL sel, struct _NSRect arg_2, char arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_832(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	char objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSSize=ff}28 */
static void 
meth_imp_833(id self, SEL sel, struct _NSRect arg_2, struct _NSSize arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_833(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	struct _NSSize objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8@12@16f36@24@28 */
static void 
meth_imp_834(id self, SEL sel, id arg_2, id arg_3, float arg_4, id arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_834(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	float objc_arg4;
	id objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8@12f36 */
static void 
meth_imp_835(id self, SEL sel, id arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_835(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8@12i16f36 */
static void 
meth_imp_836(id self, SEL sel, id arg_2, int arg_3, float arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_836(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	float objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8^{_NXStream=I**iilii^{stream_functions}^v}12i16f36 */
struct _NXStream;
static void 
meth_imp_837(id self, SEL sel, struct _NXStream  *arg_2, int arg_3, float arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NXStream=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_837(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NXStream  *objc_arg2;
	int objc_arg3;
	float objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NXStream=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8c12f36 */
static void 
meth_imp_838(id self, SEL sel, char arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_838(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8f36 */
static void 
meth_imp_839(id self, SEL sel, float arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_839(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8f36@16 */
static void 
meth_imp_840(id self, SEL sel, float arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_840(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8f36@16@20@24 */
static void 
meth_imp_841(id self, SEL sel, float arg_2, id arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_841(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8i12f36 */
static void 
meth_imp_842(id self, SEL sel, int arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_842(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8i12i16f36 */
static void 
meth_imp_843(id self, SEL sel, int arg_2, int arg_3, float arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_843(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	int objc_arg3;
	float objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8r^f12f36 */
static void 
meth_imp_844(id self, SEL sel, float  *arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_844(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float  *objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8r^f12i16f36 */
static void 
meth_imp_845(id self, SEL sel, float  *arg_2, int arg_3, float arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_845(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float  *objc_arg2;
	int objc_arg3;
	float objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8{_NSPoint=ff}12f36 */
static void 
meth_imp_846(id self, SEL sel, struct _NSPoint arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_846(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8{_NSPoint=ff}12i20f36 */
static void 
meth_imp_847(id self, SEL sel, struct _NSPoint arg_2, int arg_3, float arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_847(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	int objc_arg3;
	float objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8{_NSPoint=ff}12{_NSPoint=ff}20f36 */
static void 
meth_imp_848(id self, SEL sel, struct _NSPoint arg_2, struct _NSPoint arg_3, float arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_848(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	struct _NSPoint objc_arg3;
	float objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8{_NSPoint=ff}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}20f36 */
static void 
meth_imp_849(id self, SEL sel, struct _NSPoint arg_2, struct _NSRect arg_3, float arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_849(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	struct _NSRect objc_arg3;
	float objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v32@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12f36 */
static void 
meth_imp_850(id self, SEL sel, struct _NSRect arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_850(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8:12@16d36 */
static void 
meth_imp_851(id self, SEL sel, SEL arg_2, id arg_3, double arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_851(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	SEL objc_arg2;
	id objc_arg3;
	double objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8:12@16d36@28 */
static void 
meth_imp_852(id self, SEL sel, SEL arg_2, id arg_3, double arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_852(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	SEL objc_arg2;
	id objc_arg3;
	double objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8@12@16@20@24@28:32^v40 */
static void 
meth_imp_853(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, id arg_6, SEL arg_7, void  *arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_853(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	SEL objc_arg7;
	void  *objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8@12@16@20@24@28@32@40 */
static void 
meth_imp_854(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, id arg_6, id arg_7, id arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_854(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	id objc_arg7;
	id objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8@12@16@20@24@28@32c43 */
static void 
meth_imp_855(id self, SEL sel, id arg_2, id arg_3, id arg_4, id arg_5, id arg_6, id arg_7, char arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_855(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	id objc_arg7;
	char objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8@12I16{_NSRange=II}20i28{_NSRange=II}36 */
static void 
meth_imp_856(id self, SEL sel, id arg_2, unsigned int arg_3, struct _NSRange arg_4, int arg_5, struct _NSRange arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_856(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	unsigned int objc_arg3;
	struct _NSRange objc_arg4;
	int objc_arg5;
	struct _NSRange objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8@12^@16^c20^@24^@28^:32^I40 */
static void 
meth_imp_857(id self, SEL sel, id arg_2, id  *arg_3, char  *arg_4, id  *arg_5, id  *arg_6, SEL  *arg_7, unsigned int  *arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("^:", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_857(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id  *objc_arg3;
	char  *objc_arg4;
	id  *objc_arg5;
	id  *objc_arg6;
	SEL  *objc_arg7;
	unsigned int  *objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("^:", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8@12d36 */
static void 
meth_imp_858(id self, SEL sel, id arg_2, double arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_858(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	double objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8@12i16d36 */
static void 
meth_imp_859(id self, SEL sel, id arg_2, int arg_3, double arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_859(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	int objc_arg3;
	double objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8@12{_NSPoint=ff}16f36@28i32@40 */
static void 
meth_imp_860(id self, SEL sel, id arg_2, struct _NSPoint arg_3, float arg_4, id arg_5, int arg_6, id arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_860(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSPoint objc_arg3;
	float objc_arg4;
	id objc_arg5;
	int objc_arg6;
	id objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8@12{_NSRange=II}16I24I28^{_NSRange=II}32^I40 */
static void 
meth_imp_861(id self, SEL sel, id arg_2, struct _NSRange arg_3, unsigned int arg_4, unsigned int arg_5, struct _NSRange  *arg_6, unsigned int  *arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRange=II}", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("^I", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_861(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSRange objc_arg3;
	unsigned int objc_arg4;
	unsigned int objc_arg5;
	struct _NSRange  *objc_arg6;
	unsigned int  *objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^{_NSRange=II}", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("^I", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32c43 */
static void 
meth_imp_862(id self, SEL sel, id arg_2, struct _NSRect arg_3, id arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_862(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8@12{_NSSize=ff}16@24@28i32i40 */
static void 
meth_imp_863(id self, SEL sel, id arg_2, struct _NSSize arg_3, id arg_4, id arg_5, int arg_6, int arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_863(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSSize objc_arg3;
	id objc_arg4;
	id objc_arg5;
	int objc_arg6;
	int objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8^i12^i16^i20^i24^i28^i32@40 */
static void 
meth_imp_864(id self, SEL sel, int  *arg_2, int  *arg_3, int  *arg_4, int  *arg_5, int  *arg_6, int  *arg_7, id arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("^i", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_864(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int  *objc_arg2;
	int  *objc_arg3;
	int  *objc_arg4;
	int  *objc_arg5;
	int  *objc_arg6;
	int  *objc_arg7;
	id objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("^i", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8c12c16c20c24@28:32^v40 */
static void 
meth_imp_865(id self, SEL sel, char arg_2, char arg_3, char arg_4, char arg_5, id arg_6, SEL arg_7, void  *arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_865(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	char objc_arg3;
	char objc_arg4;
	char objc_arg5;
	id objc_arg6;
	SEL objc_arg7;
	void  *objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8c12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32@40 */
static void 
meth_imp_866(id self, SEL sel, char arg_2, struct _NSRect arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_866(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8d36 */
static void 
meth_imp_867(id self, SEL sel, double arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_867(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	double objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8d36@20 */
static void 
meth_imp_868(id self, SEL sel, double arg_2, id arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_868(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	double objc_arg2;
	id objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8d36@20:24@28 */
static void 
meth_imp_869(id self, SEL sel, double arg_2, id arg_3, SEL arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_869(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	double objc_arg2;
	id objc_arg3;
	SEL objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8d36@20:24@28@32 */
static void 
meth_imp_870(id self, SEL sel, double arg_2, id arg_3, SEL arg_4, id arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_870(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	double objc_arg2;
	id objc_arg3;
	SEL objc_arg4;
	id objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8d36c20 */
static void 
meth_imp_871(id self, SEL sel, double arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_871(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	double objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8i12i16i20{_NSRect={_NSPoint=ff}{_NSSize=ff}}28 */
static void 
meth_imp_872(id self, SEL sel, int arg_2, int arg_3, int arg_4, struct _NSRect arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_872(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	int objc_arg3;
	int objc_arg4;
	struct _NSRect objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8{_NSPoint=ff}12d36 */
static void 
meth_imp_873(id self, SEL sel, struct _NSPoint arg_2, double arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_873(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	double objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8{_NSPoint=ff}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}20i40 */
static void 
meth_imp_874(id self, SEL sel, struct _NSPoint arg_2, struct _NSRect arg_3, int arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_874(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	struct _NSRect objc_arg3;
	int objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8{_NSPoint=ff}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}20i40f36 */
static void 
meth_imp_875(id self, SEL sel, struct _NSPoint arg_2, struct _NSRect arg_3, int arg_4, float arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_875(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	struct _NSRect objc_arg3;
	int objc_arg4;
	float objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32@40 */
static void 
meth_imp_876(id self, SEL sel, struct _NSRect arg_2, id arg_3, id arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_876(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28I32@40 */
static void 
meth_imp_877(id self, SEL sel, struct _NSRect arg_2, id arg_3, unsigned int arg_4, id arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_877(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	id objc_arg3;
	unsigned int objc_arg4;
	id objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28c32i40 */
static void 
meth_imp_878(id self, SEL sel, struct _NSRect arg_2, id arg_3, char arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_878(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	id objc_arg3;
	char objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28i32i40 */
static void 
meth_imp_879(id self, SEL sel, struct _NSRect arg_2, id arg_3, int arg_4, int arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_879(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	id objc_arg3;
	int objc_arg4;
	int objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I28i32c43 */
static void 
meth_imp_880(id self, SEL sel, struct _NSRect arg_2, unsigned int arg_3, int arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_880(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	unsigned int objc_arg3;
	int objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28@32c43 */
static void 
meth_imp_881(id self, SEL sel, struct _NSRect arg_2, char arg_3, id arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_881(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	char objc_arg3;
	id objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v40@4:8@12f36f44c24 */
static void 
meth_imp_882(id self, SEL sel, id arg_2, float arg_3, float arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_882(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	float objc_arg3;
	float objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v40@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32I40@44 */
static void 
meth_imp_883(id self, SEL sel, id arg_2, struct _NSRect arg_3, id arg_4, unsigned int arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_883(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	unsigned int objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v40@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16c32@40c47 */
static void 
meth_imp_884(id self, SEL sel, id arg_2, struct _NSRect arg_3, char arg_4, id arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_884(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSRect objc_arg3;
	char objc_arg4;
	id objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v40@4:8f36f44 */
static void 
meth_imp_885(id self, SEL sel, float arg_2, float arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_885(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_arg2;
	float objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v40@4:8{_NSPoint=ff}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}20c43c47 */
static void 
meth_imp_886(id self, SEL sel, struct _NSPoint arg_2, struct _NSRect arg_3, char arg_4, char arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_886(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	struct _NSRect objc_arg3;
	char objc_arg4;
	char objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32@40@44 */
static void 
meth_imp_887(id self, SEL sel, struct _NSRect arg_2, id arg_3, id arg_4, id arg_5, id arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_887(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	id objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32 */
static void 
meth_imp_888(id self, SEL sel, struct _NSRect arg_2, struct _NSRect arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_888(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	struct _NSRect objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v44@4:8@12{_NSPoint=ff}16{_NSSize=ff}24@32@40@44c51 */
static void 
meth_imp_889(id self, SEL sel, id arg_2, struct _NSPoint arg_3, struct _NSSize arg_4, id arg_5, id arg_6, id arg_7, char arg_8)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(8);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_889(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct _NSPoint objc_arg3;
	struct _NSSize objc_arg4;
	id objc_arg5;
	id objc_arg6;
	id objc_arg7;
	char objc_arg8;
	struct objc_super super;

	if (PyTuple_Size(args) != 7) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v44@4:8d36d44 */
static void 
meth_imp_890(id self, SEL sel, double arg_2, double arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_890(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	double objc_arg2;
	double objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v44@4:8f36{_NSPoint=ff}16{_NSPoint=ff}24{_NSPoint=ff}36{_NSPoint=ff}44 */
static void 
meth_imp_891(id self, SEL sel, float arg_2, struct _NSPoint arg_3, struct _NSPoint arg_4, struct _NSPoint arg_5, struct _NSPoint arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_891(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float objc_arg2;
	struct _NSPoint objc_arg3;
	struct _NSPoint objc_arg4;
	struct _NSPoint objc_arg5;
	struct _NSPoint objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v44@4:8i12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16{_NSRect={_NSPoint=ff}{_NSSize=ff}}36 */
static void 
meth_imp_892(id self, SEL sel, int arg_2, struct _NSRect arg_3, struct _NSRect arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_892(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	struct _NSRect objc_arg3;
	struct _NSRect objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v44@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32@40i44i48 */
static void 
meth_imp_893(id self, SEL sel, struct _NSRect arg_2, id arg_3, id arg_4, id arg_5, int arg_6, int arg_7)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(7);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_893(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	id objc_arg3;
	id objc_arg4;
	id objc_arg5;
	int objc_arg6;
	int objc_arg7;
	struct objc_super super;

	if (PyTuple_Size(args) != 6) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v44@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32@48 */
static void 
meth_imp_894(id self, SEL sel, struct _NSRect arg_2, struct _NSRect arg_3, id arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_894(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	struct _NSRect objc_arg3;
	id objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v44@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32c51 */
static void 
meth_imp_895(id self, SEL sel, struct _NSRect arg_2, struct _NSRect arg_3, char arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_895(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	struct _NSRect objc_arg3;
	char objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v44@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32i48f36 */
static void 
meth_imp_896(id self, SEL sel, struct _NSRect arg_2, struct _NSRect arg_3, int arg_4, float arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_896(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	struct _NSRect objc_arg3;
	int objc_arg4;
	float objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v48@4:8@12@16{_NSPoint=ff}20{_NSSize=ff}28@40@44@48c55 */
static void 
meth_imp_897(id self, SEL sel, id arg_2, id arg_3, struct _NSPoint arg_4, struct _NSSize arg_5, id arg_6, id arg_7, id arg_8, char arg_9)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(9);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSSize=ff}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_7);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 6, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_8);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 7, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_9);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 8, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_897(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	struct _NSPoint objc_arg4;
	struct _NSSize objc_arg5;
	id objc_arg6;
	id objc_arg7;
	id objc_arg8;
	char objc_arg9;
	struct objc_super super;

	if (PyTuple_Size(args) != 8) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSSize=ff}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 5);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg7);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 6);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg8);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 7);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg9);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6, objc_arg7, objc_arg8, objc_arg9);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v48@4:8@12@16{_NSRect={_NSPoint=ff}{_NSSize=ff}}20{_NSRect={_NSPoint=ff}{_NSSize=ff}}40f36 */
static void 
meth_imp_898(id self, SEL sel, id arg_2, id arg_3, struct _NSRect arg_4, struct _NSRect arg_5, float arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_898(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	id objc_arg3;
	struct _NSRect objc_arg4;
	struct _NSRect objc_arg5;
	float objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v48@4:8i12f36f44f52 */
static void 
meth_imp_899(id self, SEL sel, int arg_2, float arg_3, float arg_4, float arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_899(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	float objc_arg3;
	float objc_arg4;
	float objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v48@4:8{_NSPoint=ff}12f36f44f52 */
static void 
meth_imp_900(id self, SEL sel, struct _NSPoint arg_2, float arg_3, float arg_4, float arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_900(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	float objc_arg3;
	float objc_arg4;
	float objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v48@4:8{_NSPoint=ff}12f36f44f52c32 */
static void 
meth_imp_901(id self, SEL sel, struct _NSPoint arg_2, float arg_3, float arg_4, float arg_5, char arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("f", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_901(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	float objc_arg3;
	float objc_arg4;
	float objc_arg5;
	char objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("f", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v48@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRange=II}28{_NSRect={_NSPoint=ff}{_NSSize=ff}}40 */
static void 
meth_imp_902(id self, SEL sel, struct _NSRect arg_2, struct _NSRange arg_3, struct _NSRect arg_4)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(4);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRange=II}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_902(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRect objc_arg2;
	struct _NSRange objc_arg3;
	struct _NSRect objc_arg4;
	struct objc_super super;

	if (PyTuple_Size(args) != 3) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRange=II}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v4@4:8 */
static void 
meth_imp_903(id self, SEL sel)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(1);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_903(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	struct objc_super super;

	if (PyTuple_Size(args) != 0) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth));
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v52@4:8i12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16{_NSRect={_NSPoint=ff}{_NSSize=ff}}36c55i56 */
static void 
meth_imp_904(id self, SEL sel, int arg_2, struct _NSRect arg_3, struct _NSRect arg_4, char arg_5, int arg_6)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(6);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_6);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 5, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_904(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	struct _NSRect objc_arg3;
	struct _NSRect objc_arg4;
	char objc_arg5;
	int objc_arg6;
	struct objc_super super;

	if (PyTuple_Size(args) != 5) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("{_NSRect={_NSPoint=ff}{_NSSize=ff}}", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 4);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg6);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5, objc_arg6);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v52@4:8{_NSPoint=ff}12d36d44d52 */
static void 
meth_imp_905(id self, SEL sel, struct _NSPoint arg_2, double arg_3, double arg_4, double arg_5)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(5);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("{_NSPoint=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_4);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 3, tmp);
	tmp = ObjC_ObjCToPython("d", &arg_5);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 4, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_905(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSPoint objc_arg2;
	double objc_arg3;
	double objc_arg4;
	double objc_arg5;
	struct objc_super super;

	if (PyTuple_Size(args) != 4) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("{_NSPoint=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 2);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg4);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 3);
	errstr = ObjC_PythonToObjC("d", v, &objc_arg5);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3, objc_arg4, objc_arg5);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v5@4:8C12 */
static void 
meth_imp_906(id self, SEL sel, unsigned char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("C", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_906(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("C", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v5@4:8c12 */
static void 
meth_imp_907(id self, SEL sel, char arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_907(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v6@4:8S12 */
static void 
meth_imp_908(id self, SEL sel, unsigned short arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_908(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned short objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8#12 */
static void 
meth_imp_909(id self, SEL sel, Class arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("#", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_909(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	Class objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("#", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8*12 */
static void 
meth_imp_910(id self, SEL sel, char* arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_910(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8:12 */
static void 
meth_imp_911(id self, SEL sel, SEL arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython(":", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_911(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	SEL objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC(":", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8@12 */
static void 
meth_imp_912(id self, SEL sel, id arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_912(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8I12 */
static void 
meth_imp_913(id self, SEL sel, unsigned int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("I", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_913(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("I", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8L12 */
static void 
meth_imp_914(id self, SEL sel, unsigned long arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("L", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_914(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned long objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("L", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^*12 */
static void 
meth_imp_915(id self, SEL sel, char*  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_915(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char*  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^@12 */
static void 
meth_imp_916(id self, SEL sel, id  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_916(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^S12 */
static void 
meth_imp_917(id self, SEL sel, unsigned short  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^S", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_917(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	unsigned short  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^S", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^f12 */
static void 
meth_imp_918(id self, SEL sel, float  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^f", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_918(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	float  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^f", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^v12 */
static void 
meth_imp_919(id self, SEL sel, void  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_919(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{?=^{_NSModalSession}c@}12 */
static void 
meth_imp_920(id self, SEL sel, struct pyobjcanonymous0  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_920(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct pyobjcanonymous0  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{?=ddd}12 */
static void 
meth_imp_921(id self, SEL sel, struct pyobjcanonymous0  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{pyobjcanonymous0=ss}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_921(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct pyobjcanonymous0  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{pyobjcanonymous0=ss}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{AEDesc=I^^{OpaqueAEDataStorageType}}12 */
static void 
meth_imp_922(id self, SEL sel, struct AEDesc  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{AEDesc=I^^{OpaqueAEDataStorageType=}}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_922(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct AEDesc  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{AEDesc=I^^{OpaqueAEDataStorageType=}}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{CGContext=}12 */
struct CGContext;
static void 
meth_imp_923(id self, SEL sel, struct CGContext  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{CGContext=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_923(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct CGContext  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{CGContext=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{FSRef=[80C]}12 */
static void 
meth_imp_924(id self, SEL sel, struct FSRef  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{FSRef=[80C]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_924(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct FSRef  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{FSRef=[80C]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{OpaqueCoreDrag=}12 */
struct OpaqueCoreDrag;
static void 
meth_imp_925(id self, SEL sel, struct OpaqueCoreDrag  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{OpaqueCoreDrag=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_925(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaqueCoreDrag  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{OpaqueCoreDrag=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{OpaqueCoreDragHandler=}12 */
struct OpaqueCoreDragHandler;
static void 
meth_imp_926(id self, SEL sel, struct OpaqueCoreDragHandler  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{OpaqueCoreDragHandler=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_926(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaqueCoreDragHandler  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{OpaqueCoreDragHandler=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{OpaqueIconRef=}12 */
struct OpaqueIconRef;
static void 
meth_imp_927(id self, SEL sel, struct OpaqueIconRef  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{OpaqueIconRef=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_927(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaqueIconRef  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{OpaqueIconRef=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{OpaqueMenuHandle=}12 */
struct OpaqueMenuHandle;
static void 
meth_imp_928(id self, SEL sel, struct OpaqueMenuHandle  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{OpaqueMenuHandle=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_928(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaqueMenuHandle  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{OpaqueMenuHandle=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{OpaquePMPageFormat=}12 */
struct OpaquePMPageFormat;
static void 
meth_imp_929(id self, SEL sel, struct OpaquePMPageFormat  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{OpaquePMPageFormat=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_929(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaquePMPageFormat  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{OpaquePMPageFormat=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{OpaquePMPrintSettings=}12 */
struct OpaquePMPrintSettings;
static void 
meth_imp_930(id self, SEL sel, struct OpaquePMPrintSettings  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{OpaquePMPrintSettings=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_930(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct OpaquePMPrintSettings  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{OpaquePMPrintSettings=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}12 */
struct _NSModalSession;
static void 
meth_imp_931(id self, SEL sel, struct _NSModalSession  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSModalSession=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_931(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSModalSession  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSModalSession=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{_NSRefCountedRunArray=IIIIII[0{_NSRunArrayItem=I@}]}12 */
static void 
meth_imp_932(id self, SEL sel, struct _NSRefCountedRunArray  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSRefCountedRunArray=IIIIII[0{_NSRunArrayItem=I@}]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_932(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSRefCountedRunArray  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSRefCountedRunArray=IIIIII[0{_NSRunArrayItem=I@}]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{_NSSortState=iIIII[4@]}12 */
static void 
meth_imp_933(id self, SEL sel, struct _NSSortState  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSSortState=iIIII[4@]}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_933(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSSortState  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSSortState=iIIII[4@]}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{_NSZone=}12 */
struct _NSZone;
static void 
meth_imp_934(id self, SEL sel, struct _NSZone  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSZone=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_934(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSZone  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSZone=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{__CFHTTPMessage=}12 */
struct __CFHTTPMessage;
static void 
meth_imp_935(id self, SEL sel, struct __CFHTTPMessage  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{__CFHTTPMessage=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_935(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFHTTPMessage  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{__CFHTTPMessage=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{__CFString=}12 */
struct __CFString;
static void 
meth_imp_936(id self, SEL sel, struct __CFString  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{__CFString=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_936(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct __CFString  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{__CFString=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8^{tiff=*^{_NXStream}sccsll{?=IIIIIISSSSSSSSSSIIIffSSffII[2S]ISSSSI^S^S^S^S[3^S]*********[2I]II^I^I[2S]^f[2S]S^f^f^f[4^S]S[2S]**I^v}{?=SSL}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}12 */
static void 
meth_imp_937(id self, SEL sel, struct tiff  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{tiff=*^{_NXStream=}sccsll{pyobjcanonymous0=ss}{pyobjcanonymous0=ss}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_937(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct tiff  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{tiff=*^{_NXStream=}sccsll{pyobjcanonymous0=ss}{pyobjcanonymous0=ss}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8i12 */
static void 
meth_imp_938(id self, SEL sel, int arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_938(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8l12 */
static void 
meth_imp_939(id self, SEL sel, long arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("l", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_939(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	long objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("l", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8r*12 */
static void 
meth_imp_940(id self, SEL sel, char* arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("*", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_940(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char* objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("*", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v8@4:8r^v12 */
static void 
meth_imp_941(id self, SEL sel, void  *arg_2)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(2);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^v", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_941(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	void  *objc_arg2;
	struct objc_super super;

	if (PyTuple_Size(args) != 1) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^v", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v9@4:8@12c16 */
static void 
meth_imp_942(id self, SEL sel, id arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("@", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_942(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	id objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("@", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v9@4:8^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}12c16 */
struct _NSModalSession;
static void 
meth_imp_943(id self, SEL sel, struct _NSModalSession  *arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSModalSession=}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_943(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSModalSession  *objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSModalSession=}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v9@4:8^{_NSSize=ff}12c16 */
static void 
meth_imp_944(id self, SEL sel, struct _NSSize  *arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("^{_NSSize=ff}", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_944(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	struct _NSSize  *objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("^{_NSSize=ff}", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v9@4:8c12c16 */
static void 
meth_imp_945(id self, SEL sel, char arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_945(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	char objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


/* signature: v9@4:8i12c16 */
static void 
meth_imp_946(id self, SEL sel, int arg_2, char arg_3)
{
	PyObject* arglist;
	PyObject* retval;
	PyObject* tmp;

	arglist = PyTuple_New(3);
	if (arglist == NULL) ObjCErr_ToObjC();

	tmp = ObjC_ObjCToPython("@", &self);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 0, tmp);
	tmp = ObjC_ObjCToPython("i", &arg_2);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 1, tmp);
	tmp = ObjC_ObjCToPython("c", &arg_3);
	if (tmp == NULL) ObjCErr_ToObjC();
	PyTuple_SetItem(arglist, 2, tmp);

	retval = ObjC_CallPython(self, sel, arglist);
	Py_DECREF(arglist);
	if (retval == NULL) ObjCErr_ToObjC();
}
static PyObject* super_946(PyObject* meth, PyObject* self, PyObject* args)
{
	id objc_self;
	const char* errstr;
	PyObject* v;
	int objc_arg2;
	char objc_arg3;
	struct objc_super super;

	if (PyTuple_Size(args) != 2) {
		PyErr_SetString(PyExc_TypeError, "Wrong argcount");
		return NULL;
	}
	errstr = ObjC_PythonToObjC("@", self, &objc_self);
	if (errstr != NULL) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert self");
		return NULL;
	} 	super.receiver = objc_self;
	super.class = ObjCSelector_GetClass(meth);
	v = PyTuple_GetItem(args, 0);
	errstr = ObjC_PythonToObjC("i", v, &objc_arg2);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	v = PyTuple_GetItem(args, 1);
	errstr = ObjC_PythonToObjC("c", v, &objc_arg3);
	if (errstr) {
		PyErr_SetString(PyExc_TypeError, "Cannot convert argument");
	return NULL;
	}
	NS_DURING
		(void)objc_msgSendSuper(&super, ObjCSelector_GetSelector(meth), objc_arg2, objc_arg3);
	NS_HANDLER
		ObjCErr_FromObjC(localException);
	NS_ENDHANDLER
	if (PyErr_Occurred()) return NULL;
	Py_INCREF(Py_None);
	return Py_None;
}


static struct method_table {
	char* signature;
	superfunc call_super;
	IMP implementation;
} method_table[] = {
	{ "#12@4:8@12@16", (superfunc)super_0, (IMP)meth_imp_0 },
	{ "#4@4:8", (superfunc)super_1, (IMP)meth_imp_1 },
	{ "#8@4:8@12", (superfunc)super_2, (IMP)meth_imp_2 },
	{ "#8@4:8I12", (superfunc)super_3, (IMP)meth_imp_3 },
	{ "*12@4:8@12^I16", (superfunc)super_4, (IMP)meth_imp_4 },
	{ "*4@4:8", (superfunc)super_5, (IMP)meth_imp_5 },
	{ "*8@4:8r*12", (superfunc)super_6, (IMP)meth_imp_6 },
	{ ":4@4:8", (superfunc)super_7, (IMP)meth_imp_7 },
	{ ":8@4:8@12", (superfunc)super_8, (IMP)meth_imp_8 },
	{ "@10@4:8S12S16", (superfunc)super_9, (IMP)meth_imp_9 },
	{ "@120@4:8{_CGSEventRecord=SSII{CGPoint=ff}{CGPoint=ff}QI^v^v(?={?=CCsiCcCCss(?={_CGSTabletPointData=iiiSS{?=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})[4i]}{?=CCsiCcCCss(?={_CGSTabletPointData=iiiSS{?=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})[4i]}{?=ssSSSsssI[11i]}{?=ssii[13i]}{?=SSIIi[12i]}{?=ssssi[13i]}{?=iiiSS{?=ss}SsSsss[8i]}{?=SSSSSSIQICCs[8i]}{?=ss(?=[15f][15i][30s][60c])})}16", (superfunc)super_10, (IMP)meth_imp_10 },
	{ "@124@4:8{_CGSEventRecord=SSII{CGPoint=ff}{CGPoint=ff}QI^v^v(?={?=CCsiCcCCss(?={_CGSTabletPointData=iiiSS{?=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})[4i]}{?=CCsiCcCCss(?={_CGSTabletPointData=iiiSS{?=ss}SsSsss}{_CGSTabletProximityData=SSSSSSIQICCs})[4i]}{?=ssSSSsssI[11i]}{?=ssii[13i]}{?=SSIIi[12i]}{?=ssssi[13i]}{?=iiiSS{?=ss}SsSsss[8i]}{?=SSSSSSIQICCs[8i]}{?=ss(?=[15f][15i][30s][60c])})}16^v128", (superfunc)super_11, (IMP)meth_imp_11 },
	{ "@12@4:8*12I16", (superfunc)super_12, (IMP)meth_imp_12 },
	{ "@12@4:8*12i16", (superfunc)super_13, (IMP)meth_imp_13 },
	{ "@12@4:8*16", (superfunc)super_14, (IMP)meth_imp_14 },
	{ "@12@4:8:12@16", (superfunc)super_15, (IMP)meth_imp_15 },
	{ "@12@4:8:12^:16", (superfunc)super_16, (IMP)meth_imp_16 },
	{ "@12@4:8:12^v16", (superfunc)super_17, (IMP)meth_imp_17 },
	{ "@12@4:8@12#16", (superfunc)super_18, (IMP)meth_imp_18 },
	{ "@12@4:8@12*16", (superfunc)super_19, (IMP)meth_imp_19 },
	{ "@12@4:8@12@16", (superfunc)super_20, (IMP)meth_imp_20 },
	{ "@12@4:8@12I16", (superfunc)super_21, (IMP)meth_imp_21 },
	{ "@12@4:8@12^{?=^SI^SI^SI}16", (superfunc)super_22, (IMP)meth_imp_22 },
	{ "@12@4:8@12^{_NSZone=}16", (superfunc)super_23, (IMP)meth_imp_23 },
	{ "@12@4:8@12i16", (superfunc)super_24, (IMP)meth_imp_24 },
	{ "@12@4:8@12r^f16", (superfunc)super_25, (IMP)meth_imp_25 },
	{ "@12@4:8@12r^{FSRef=[80C]}16", (superfunc)super_26, (IMP)meth_imp_26 },
	{ "@12@4:8@12r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_27, (IMP)meth_imp_27 },
	{ "@12@4:8@16", (superfunc)super_28, (IMP)meth_imp_28 },
	{ "@12@4:8I12:16", (superfunc)super_29, (IMP)meth_imp_29 },
	{ "@12@4:8I12@16", (superfunc)super_30, (IMP)meth_imp_30 },
	{ "@12@4:8I12I16", (superfunc)super_31, (IMP)meth_imp_31 },
	{ "@12@4:8I12^I16", (superfunc)super_32, (IMP)meth_imp_32 },
	{ "@12@4:8I12^{_NSRange=II}16", (superfunc)super_33, (IMP)meth_imp_33 },
	{ "@12@4:8L12L16", (superfunc)super_34, (IMP)meth_imp_34 },
	{ "@12@4:8Q12", (superfunc)super_35, (IMP)meth_imp_35 },
	{ "@12@4:8S12@16", (superfunc)super_36, (IMP)meth_imp_36 },
	{ "@12@4:8S12i16", (superfunc)super_37, (IMP)meth_imp_37 },
	{ "@12@4:8^?12^v16", (superfunc)super_38, (IMP)meth_imp_38 },
	{ "@12@4:8^?12i16", (superfunc)super_39, (IMP)meth_imp_39 },
	{ "@12@4:8^@12@16", (superfunc)super_40, (IMP)meth_imp_40 },
	{ "@12@4:8^@12I16", (superfunc)super_41, (IMP)meth_imp_41 },
	{ "@12@4:8^S12I16", (superfunc)super_42, (IMP)meth_imp_42 },
	{ "@12@4:8^i12^i16", (superfunc)super_43, (IMP)meth_imp_43 },
	{ "@12@4:8^v12I16", (superfunc)super_44, (IMP)meth_imp_44 },
	{ "@12@4:8^{FSRef=[80C]}12i16", (superfunc)super_45, (IMP)meth_imp_45 },
	{ "@12@4:8^{_ProtocolTemplate=#*^{objc_protocol_list}^{objc_method_description_list}^{objc_method_description_list}}12i16", (superfunc)super_46, (IMP)meth_imp_46 },
	{ "@12@4:8^{hostent=*^*ii^*}12@16", (superfunc)super_47, (IMP)meth_imp_47 },
	{ "@12@4:8c12@16", (superfunc)super_48, (IMP)meth_imp_48 },
	{ "@12@4:8c12i16", (superfunc)super_49, (IMP)meth_imp_49 },
	{ "@12@4:8i12@16", (superfunc)super_50, (IMP)meth_imp_50 },
	{ "@12@4:8i12i16", (superfunc)super_51, (IMP)meth_imp_51 },
	{ "@12@4:8i12r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_52, (IMP)meth_imp_52 },
	{ "@12@4:8q12", (superfunc)super_53, (IMP)meth_imp_53 },
	{ "@12@4:8r*12I16", (superfunc)super_54, (IMP)meth_imp_54 },
	{ "@12@4:8r*16", (superfunc)super_55, (IMP)meth_imp_55 },
	{ "@12@4:8r^S12I16", (superfunc)super_56, (IMP)meth_imp_56 },
	{ "@12@4:8r^v12I16", (superfunc)super_57, (IMP)meth_imp_57 },
	{ "@12@4:8r^v12r*16", (superfunc)super_58, (IMP)meth_imp_58 },
	{ "@12@4:8r^{_NSSize=ff}12@16", (superfunc)super_59, (IMP)meth_imp_59 },
	{ "@12@4:8s12@16", (superfunc)super_60, (IMP)meth_imp_60 },
	{ "@12@4:8{CGPoint=ff}12", (superfunc)super_61, (IMP)meth_imp_61 },
	{ "@12@4:8{NSButtonState=iccc}12", (superfunc)super_62, (IMP)meth_imp_62 },
	{ "@12@4:8{_NSPoint=ff}12", (superfunc)super_63, (IMP)meth_imp_63 },
	{ "@12@4:8{_NSRange=II}12", (superfunc)super_64, (IMP)meth_imp_64 },
	{ "@12@4:8{_NSSize=ff}12", (superfunc)super_65, (IMP)meth_imp_65 },
	{ "@13@4:8*12I16c20", (superfunc)super_66, (IMP)meth_imp_66 },
	{ "@13@4:8@12@16c20", (superfunc)super_67, (IMP)meth_imp_67 },
	{ "@13@4:8@12^I16c20", (superfunc)super_68, (IMP)meth_imp_68 },
	{ "@13@4:8@12^{?=^SI^SI^SI}16c20", (superfunc)super_69, (IMP)meth_imp_69 },
	{ "@13@4:8@12c16c20", (superfunc)super_70, (IMP)meth_imp_70 },
	{ "@13@4:8^@12c16c20", (superfunc)super_71, (IMP)meth_imp_71 },
	{ "@13@4:8^S12I16c20", (superfunc)super_72, (IMP)meth_imp_72 },
	{ "@13@4:8^{FSRef=[80C]}12c16c20", (superfunc)super_73, (IMP)meth_imp_73 },
	{ "@13@4:8i12i16c20", (superfunc)super_74, (IMP)meth_imp_74 },
	{ "@13@4:8r^v12I16c20", (superfunc)super_75, (IMP)meth_imp_75 },
	{ "@13@4:8{_NSPoint=ff}12c20", (superfunc)super_76, (IMP)meth_imp_76 },
	{ "@13@4:8{_NSRange=II}12c20", (superfunc)super_77, (IMP)meth_imp_77 },
	{ "@14@4:8@12@16S20", (superfunc)super_78, (IMP)meth_imp_78 },
	{ "@14@4:8@12^{tiff=*^{_NXStream}sccsll{?=IIIIIISSSSSSSSSSIIIffSSffII[2S]ISSSSI^S^S^S^S[3^S]*********[2I]II^I^I[2S]^f[2S]S^f^f^f[4^S]S[2S]**I^v}{?=SSL}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}16s20", (superfunc)super_79, (IMP)meth_imp_79 },
	{ "@16@4:8*12*20", (superfunc)super_80, (IMP)meth_imp_80 },
	{ "@16@4:8:12@16@20", (superfunc)super_81, (IMP)meth_imp_81 },
	{ "@16@4:8@12:16@20", (superfunc)super_82, (IMP)meth_imp_82 },
	{ "@16@4:8@12@16*20", (superfunc)super_83, (IMP)meth_imp_83 },
	{ "@16@4:8@12@16@20", (superfunc)super_84, (IMP)meth_imp_84 },
	{ "@16@4:8@12@16I20", (superfunc)super_85, (IMP)meth_imp_85 },
	{ "@16@4:8@12@16^c20", (superfunc)super_86, (IMP)meth_imp_86 },
	{ "@16@4:8@12@16^{_NSPoint=ff}20", (superfunc)super_87, (IMP)meth_imp_87 },
	{ "@16@4:8@12@16^{_NSZone=}20", (superfunc)super_88, (IMP)meth_imp_88 },
	{ "@16@4:8@12@16i20", (superfunc)super_89, (IMP)meth_imp_89 },
	{ "@16@4:8@12@20", (superfunc)super_90, (IMP)meth_imp_90 },
	{ "@16@4:8@12I16@20", (superfunc)super_91, (IMP)meth_imp_91 },
	{ "@16@4:8@12I16I20", (superfunc)super_92, (IMP)meth_imp_92 },
	{ "@16@4:8@12I16^{_NSRange=II}20", (superfunc)super_93, (IMP)meth_imp_93 },
	{ "@16@4:8@12I16i20", (superfunc)super_94, (IMP)meth_imp_94 },
	{ "@16@4:8@12^@16^{_NSZone=}20", (superfunc)super_95, (IMP)meth_imp_95 },
	{ "@16@4:8@12^{OpaquePMPageFormat=}16^{OpaquePMPrintSettings=}20", (superfunc)super_96, (IMP)meth_imp_96 },
	{ "@16@4:8@12i16:20", (superfunc)super_97, (IMP)meth_imp_97 },
	{ "@16@4:8@12i16@20", (superfunc)super_98, (IMP)meth_imp_98 },
	{ "@16@4:8@12i16I20", (superfunc)super_99, (IMP)meth_imp_99 },
	{ "@16@4:8@12i16i20", (superfunc)super_100, (IMP)meth_imp_100 },
	{ "@16@4:8@12i16r*20", (superfunc)super_101, (IMP)meth_imp_101 },
	{ "@16@4:8@12r*16I20", (superfunc)super_102, (IMP)meth_imp_102 },
	{ "@16@4:8@12{_NSPoint=ff}16", (superfunc)super_103, (IMP)meth_imp_103 },
	{ "@16@4:8@12{_NSRange=II}16", (superfunc)super_104, (IMP)meth_imp_104 },
	{ "@16@4:8I12^{_NSRange=II}16^I20", (superfunc)super_105, (IMP)meth_imp_105 },
	{ "@16@4:8I12r^v16L20", (superfunc)super_106, (IMP)meth_imp_106 },
	{ "@16@4:8I12{_NSRange=II}16", (superfunc)super_107, (IMP)meth_imp_107 },
	{ "@16@4:8S12I16@20", (superfunc)super_108, (IMP)meth_imp_108 },
	{ "@16@4:8S12S16@20", (superfunc)super_109, (IMP)meth_imp_109 },
	{ "@16@4:8^?12^?16:20", (superfunc)super_110, (IMP)meth_imp_110 },
	{ "@16@4:8^?12^?16I20", (superfunc)super_111, (IMP)meth_imp_111 },
	{ "@16@4:8^?12^v16@20", (superfunc)super_112, (IMP)meth_imp_112 },
	{ "@16@4:8^@12^@16I20", (superfunc)super_113, (IMP)meth_imp_113 },
	{ "@16@4:8^@12^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}20", (superfunc)super_114, (IMP)meth_imp_114 },
	{ "@16@4:8^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12r*16*20", (superfunc)super_115, (IMP)meth_imp_115 },
	{ "@16@4:8^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12r*16r*20", (superfunc)super_116, (IMP)meth_imp_116 },
	{ "@16@4:8i12@16^i20", (superfunc)super_117, (IMP)meth_imp_117 },
	{ "@16@4:8i12@16i20", (superfunc)super_118, (IMP)meth_imp_118 },
	{ "@16@4:8i12i16@20", (superfunc)super_119, (IMP)meth_imp_119 },
	{ "@16@4:8i12i16i20", (superfunc)super_120, (IMP)meth_imp_120 },
	{ "@16@4:8i12r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16I20", (superfunc)super_121, (IMP)meth_imp_121 },
	{ "@16@4:8i12{_NSRange=II}16", (superfunc)super_122, (IMP)meth_imp_122 },
	{ "@16@4:8r*12I16I20", (superfunc)super_123, (IMP)meth_imp_123 },
	{ "@16@4:8{_NSRange=II}12^{_NSZone=}20", (superfunc)super_124, (IMP)meth_imp_124 },
	{ "@16@4:8{_NSSize=ff}12@20", (superfunc)super_125, (IMP)meth_imp_125 },
	{ "@16@4:8{_NSSize=ff}12i20", (superfunc)super_126, (IMP)meth_imp_126 },
	{ "@17@4:8@12@16@20c24", (superfunc)super_127, (IMP)meth_imp_127 },
	{ "@17@4:8@12@16i20c24", (superfunc)super_128, (IMP)meth_imp_128 },
	{ "@17@4:8@12^I16I20c24", (superfunc)super_129, (IMP)meth_imp_129 },
	{ "@17@4:8I12@16@20c24", (superfunc)super_130, (IMP)meth_imp_130 },
	{ "@17@4:8Q12s20c24", (superfunc)super_131, (IMP)meth_imp_131 },
	{ "@17@4:8^{FSCatalogInfo=SsIICCCC{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}{UTCDateTime=SIS}[4I][16C][16C]QQQQII}12@16^{FSRef=[80C]}20c24", (superfunc)super_132, (IMP)meth_imp_132 },
	{ "@17@4:8^{_SelectionAnchor=iii}12^{_SelectionAnchor=iii}16c20c24", (superfunc)super_133, (IMP)meth_imp_133 },
	{ "@17@4:8c12i16i20c24", (superfunc)super_134, (IMP)meth_imp_134 },
	{ "@20@4:8#12@16@20:24", (superfunc)super_135, (IMP)meth_imp_135 },
	{ "@20@4:8:12i16@20@24", (superfunc)super_136, (IMP)meth_imp_136 },
	{ "@20@4:8@12:16@20i24", (superfunc)super_137, (IMP)meth_imp_137 },
	{ "@20@4:8@12@16:20@24", (superfunc)super_138, (IMP)meth_imp_138 },
	{ "@20@4:8@12@16@20@24", (superfunc)super_139, (IMP)meth_imp_139 },
	{ "@20@4:8@12@16@20^@24", (superfunc)super_140, (IMP)meth_imp_140 },
	{ "@20@4:8@12@16@20^{_NSZone=}24", (superfunc)super_141, (IMP)meth_imp_141 },
	{ "@20@4:8@12@16@20i24", (superfunc)super_142, (IMP)meth_imp_142 },
	{ "@20@4:8@12@16I20@24", (superfunc)super_143, (IMP)meth_imp_143 },
	{ "@20@4:8@12@16c20@24", (superfunc)super_144, (IMP)meth_imp_144 },
	{ "@20@4:8@12@16i20i24", (superfunc)super_145, (IMP)meth_imp_145 },
	{ "@20@4:8@12i16i20@24", (superfunc)super_146, (IMP)meth_imp_146 },
	{ "@20@4:8@12{_NSRange=II}16i24", (superfunc)super_147, (IMP)meth_imp_147 },
	{ "@20@4:8I12@16@20^{_NSZone=}24", (superfunc)super_148, (IMP)meth_imp_148 },
	{ "@20@4:8I12^{_NSRange=II}16{_NSRange=II}20", (superfunc)super_149, (IMP)meth_imp_149 },
	{ "@20@4:8^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12r*16^*20i24", (superfunc)super_150, (IMP)meth_imp_150 },
	{ "@20@4:8^{__CFSocket=}12i16i20i24", (superfunc)super_151, (IMP)meth_imp_151 },
	{ "@20@4:8i12i16i20@24", (superfunc)super_152, (IMP)meth_imp_152 },
	{ "@20@4:8i12i16i20i24", (superfunc)super_153, (IMP)meth_imp_153 },
	{ "@20@4:8r*12r*16r*20^{?=b4b1b24(?=*^{?}^{__CFDictionary})}24", (superfunc)super_154, (IMP)meth_imp_154 },
	{ "@20@4:8{_NSRange=II}12@20@24", (superfunc)super_155, (IMP)meth_imp_155 },
	{ "@20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12", (superfunc)super_156, (IMP)meth_imp_156 },
	{ "@21@4:8@12@16@20@24c28", (superfunc)super_157, (IMP)meth_imp_157 },
	{ "@21@4:8^@12I16@20c24c28", (superfunc)super_158, (IMP)meth_imp_158 },
	{ "@21@4:8^v12I16c20c24c28", (superfunc)super_159, (IMP)meth_imp_159 },
	{ "@21@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28", (superfunc)super_160, (IMP)meth_imp_160 },
	{ "@21@4:8{_NSSize=ff}12i20c24c28", (superfunc)super_161, (IMP)meth_imp_161 },
	{ "@22@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12s28", (superfunc)super_162, (IMP)meth_imp_162 },
	{ "@24@4:8*12*16*20*24*28", (superfunc)super_163, (IMP)meth_imp_163 },
	{ "@24@4:8@12@16@20@24@28", (superfunc)super_164, (IMP)meth_imp_164 },
	{ "@24@4:8@12@16@20i24@28", (superfunc)super_165, (IMP)meth_imp_165 },
	{ "@24@4:8@12@16@20{_NSPoint=ff}24", (superfunc)super_166, (IMP)meth_imp_166 },
	{ "@24@4:8@12@16I20@24@28", (superfunc)super_167, (IMP)meth_imp_167 },
	{ "@24@4:8@12@16{_NSRange=II}20@28", (superfunc)super_168, (IMP)meth_imp_168 },
	{ "@24@4:8@12I16^{_NSRange=II}20{_NSRange=II}24", (superfunc)super_169, (IMP)meth_imp_169 },
	{ "@24@4:8@12i16{_NSPoint=ff}20^v28", (superfunc)super_170, (IMP)meth_imp_170 },
	{ "@24@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_171, (IMP)meth_imp_171 },
	{ "@24@4:8I12I16@20s24i28", (superfunc)super_172, (IMP)meth_imp_172 },
	{ "@24@4:8^v12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_173, (IMP)meth_imp_173 },
	{ "@24@4:8i12@16@20@24i28", (superfunc)super_174, (IMP)meth_imp_174 },
	{ "@24@4:8i12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_175, (IMP)meth_imp_175 },
	{ "@24@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I16i20c24@28", (superfunc)super_176, (IMP)meth_imp_176 },
	{ "@24@4:8{?=b8b4b1b1b18[8S]}12", (superfunc)super_177, (IMP)meth_imp_177 },
	{ "@24@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28", (superfunc)super_178, (IMP)meth_imp_178 },
	{ "@24@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12i28", (superfunc)super_179, (IMP)meth_imp_179 },
	{ "@25@4:8*12*16*20*24*28c32", (superfunc)super_180, (IMP)meth_imp_180 },
	{ "@25@4:8@12@16@20@24^@28c32", (superfunc)super_181, (IMP)meth_imp_181 },
	{ "@25@4:8@12@16i20i24^{_SelectionAnchor=iii}28c32", (superfunc)super_182, (IMP)meth_imp_182 },
	{ "@25@4:8i12s16c20c24c28c32", (superfunc)super_183, (IMP)meth_imp_183 },
	{ "@25@4:8{_NSSize=ff}12i20c24c28c32", (superfunc)super_184, (IMP)meth_imp_184 },
	{ "@28@4:8@12@16@20@24@28@32", (superfunc)super_185, (IMP)meth_imp_185 },
	{ "@28@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32", (superfunc)super_186, (IMP)meth_imp_186 },
	{ "@28@4:8i12i16i20i24i28i32", (superfunc)super_187, (IMP)meth_imp_187 },
	{ "@28@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I16i20c24@28@32", (superfunc)super_188, (IMP)meth_imp_188 },
	{ "@28@4:8{_NSRange=II}12@20@24{_NSRange=II}28", (superfunc)super_189, (IMP)meth_imp_189 },
	{ "@28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32", (superfunc)super_190, (IMP)meth_imp_190 },
	{ "@28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28i32", (superfunc)super_191, (IMP)meth_imp_191 },
	{ "@28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I28@32", (superfunc)super_192, (IMP)meth_imp_192 },
	{ "@32@4:8@12@16f36", (superfunc)super_193, (IMP)meth_imp_193 },
	{ "@32@4:8@12I16i20f36", (superfunc)super_194, (IMP)meth_imp_194 },
	{ "@32@4:8@12f36", (superfunc)super_195, (IMP)meth_imp_195 },
	{ "@32@4:8@12f36@20{_NSPoint=ff}24", (superfunc)super_196, (IMP)meth_imp_196 },
	{ "@32@4:8@12f36r^f20", (superfunc)super_197, (IMP)meth_imp_197 },
	{ "@32@4:8@12f36r^f20I24", (superfunc)super_198, (IMP)meth_imp_198 },
	{ "@32@4:8@12f36r^f20i24", (superfunc)super_199, (IMP)meth_imp_199 },
	{ "@32@4:8@12i16f36", (superfunc)super_200, (IMP)meth_imp_200 },
	{ "@32@4:8^{?=*i}12^*16^*20f36", (superfunc)super_201, (IMP)meth_imp_201 },
	{ "@32@4:8f36", (superfunc)super_202, (IMP)meth_imp_202 },
	{ "@32@4:8f36@16", (superfunc)super_203, (IMP)meth_imp_203 },
	{ "@32@4:8i12f36", (superfunc)super_204, (IMP)meth_imp_204 },
	{ "@32@4:8i12f36r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}20r^{_NSPoint=ff}24", (superfunc)super_205, (IMP)meth_imp_205 },
	{ "@36@4:8@12:16@20@24@28@32I40", (superfunc)super_206, (IMP)meth_imp_206 },
	{ "@36@4:8@12@16c20@24@28:32I40", (superfunc)super_207, (IMP)meth_imp_207 },
	{ "@36@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32@40", (superfunc)super_208, (IMP)meth_imp_208 },
	{ "@36@4:8d36", (superfunc)super_209, (IMP)meth_imp_209 },
	{ "@36@4:8d36@20", (superfunc)super_210, (IMP)meth_imp_210 },
	{ "@36@4:8d36@20:24@28c32", (superfunc)super_211, (IMP)meth_imp_211 },
	{ "@36@4:8d36@20c24", (superfunc)super_212, (IMP)meth_imp_212 },
	{ "@36@4:8i12@16@20@24@28@32*40", (superfunc)super_213, (IMP)meth_imp_213 },
	{ "@36@4:8i12I16I20I24I28I32@40", (superfunc)super_214, (IMP)meth_imp_214 },
	{ "@36@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@16@20@24@28i32i40", (superfunc)super_215, (IMP)meth_imp_215 },
	{ "@36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28I32@40", (superfunc)super_216, (IMP)meth_imp_216 },
	{ "@36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I28i32c43", (superfunc)super_217, (IMP)meth_imp_217 },
	{ "@40@4:8@12d36@24:28@32c43c47", (superfunc)super_218, (IMP)meth_imp_218 },
	{ "@40@4:8@12{_NSSize=ff}16f36f44{_NSPoint=ff}36", (superfunc)super_219, (IMP)meth_imp_219 },
	{ "@40@4:8f36f44", (superfunc)super_220, (IMP)meth_imp_220 },
	{ "@40@4:8f36f44c20", (superfunc)super_221, (IMP)meth_imp_221 },
	{ "@40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I28i32c43@44", (superfunc)super_222, (IMP)meth_imp_222 },
	{ "@40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12i28#32i40i44", (superfunc)super_223, (IMP)meth_imp_223 },
	{ "@40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12i28@32i40i44", (superfunc)super_224, (IMP)meth_imp_224 },
	{ "@48@4:8^*12i16i20i24i28c32c43@44i48i52", (superfunc)super_225, (IMP)meth_imp_225 },
	{ "@48@4:8i12{_NSPoint=ff}16I24d36i40@44i48i52f44", (superfunc)super_226, (IMP)meth_imp_226 },
	{ "@4@4:8", (superfunc)super_227, (IMP)meth_imp_227 },
	{ "@52@4:8i12{_NSPoint=ff}16I24d36i40@44i48i52^v56", (superfunc)super_228, (IMP)meth_imp_228 },
	{ "@52@4:8i12{_NSPoint=ff}16I24d36i40@44s50i52i56", (superfunc)super_229, (IMP)meth_imp_229 },
	{ "@56@4:8^*12i16i20i24i28c32c43@44i48i52{_NSSize=ff}56", (superfunc)super_230, (IMP)meth_imp_230 },
	{ "@56@4:8f36f44f52f60", (superfunc)super_231, (IMP)meth_imp_231 },
	{ "@56@4:8i12{_NSPoint=ff}16I24d36i40@44@48@52c59S62", (superfunc)super_232, (IMP)meth_imp_232 },
	{ "@5@4:8C12", (superfunc)super_233, (IMP)meth_imp_233 },
	{ "@5@4:8c12", (superfunc)super_234, (IMP)meth_imp_234 },
	{ "@64@4:8f36f44f52f60f68", (superfunc)super_235, (IMP)meth_imp_235 },
	{ "@6@4:8S12", (superfunc)super_236, (IMP)meth_imp_236 },
	{ "@6@4:8s12", (superfunc)super_237, (IMP)meth_imp_237 },
	{ "@8@4:8#12", (superfunc)super_238, (IMP)meth_imp_238 },
	{ "@8@4:8*12", (superfunc)super_239, (IMP)meth_imp_239 },
	{ "@8@4:8:12", (superfunc)super_240, (IMP)meth_imp_240 },
	{ "@8@4:8@12", (superfunc)super_241, (IMP)meth_imp_241 },
	{ "@8@4:8I12", (superfunc)super_242, (IMP)meth_imp_242 },
	{ "@8@4:8L12", (superfunc)super_243, (IMP)meth_imp_243 },
	{ "@8@4:8^c12", (superfunc)super_244, (IMP)meth_imp_244 },
	{ "@8@4:8^i12", (superfunc)super_245, (IMP)meth_imp_245 },
	{ "@8@4:8^v12", (superfunc)super_246, (IMP)meth_imp_246 },
	{ "@8@4:8^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12", (superfunc)super_247, (IMP)meth_imp_247 },
	{ "@8@4:8^{FSRef=[80C]}12", (superfunc)super_248, (IMP)meth_imp_248 },
	{ "@8@4:8^{NSCharSetPrivateStruct=i[4i]iiii[1i]}12", (superfunc)super_249, (IMP)meth_imp_249 },
	{ "@8@4:8^{_NSPoint=ff}12", (superfunc)super_250, (IMP)meth_imp_250 },
	{ "@8@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12", (superfunc)super_251, (IMP)meth_imp_251 },
	{ "@8@4:8^{_NSRefCountedRunArray=IIIIII[0{_NSRunArrayItem=I@}]}12", (superfunc)super_252, (IMP)meth_imp_252 },
	{ "@8@4:8^{_NSRulebookSetHeader=i[4L]iiii[1i]}12", (superfunc)super_253, (IMP)meth_imp_253 },
	{ "@8@4:8^{_NSSize=ff}12", (superfunc)super_254, (IMP)meth_imp_254 },
	{ "@8@4:8^{_NSStringBuffer=II@II[32S]S}12", (superfunc)super_255, (IMP)meth_imp_255 },
	{ "@8@4:8^{_NSZone=}12", (superfunc)super_256, (IMP)meth_imp_256 },
	{ "@8@4:8^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}12", (superfunc)super_257, (IMP)meth_imp_257 },
	{ "@8@4:8^{__CFNotificationCenter=}12", (superfunc)super_258, (IMP)meth_imp_258 },
	{ "@8@4:8^{_object=i^{_typeobject}}12", (superfunc)super_259, (IMP)meth_imp_259 },
	{ "@8@4:8^{hostent=*^*ii^*}12", (superfunc)super_260, (IMP)meth_imp_260 },
	{ "@8@4:8^{stat=iISSIIi{timespec=ii}{timespec=ii}{timespec=ii}qqIIIi[2q]}12", (superfunc)super_261, (IMP)meth_imp_261 },
	{ "@8@4:8i12", (superfunc)super_262, (IMP)meth_imp_262 },
	{ "@8@4:8l12", (superfunc)super_263, (IMP)meth_imp_263 },
	{ "@8@4:8r*12", (superfunc)super_264, (IMP)meth_imp_264 },
	{ "@8@4:8r^v12", (superfunc)super_265, (IMP)meth_imp_265 },
	{ "@8@4:8r^{FSRef=[80C]}12", (superfunc)super_266, (IMP)meth_imp_266 },
	{ "@8@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12", (superfunc)super_267, (IMP)meth_imp_267 },
	{ "@9@4:8:12c16", (superfunc)super_268, (IMP)meth_imp_268 },
	{ "@9@4:8@12c16", (superfunc)super_269, (IMP)meth_imp_269 },
	{ "@9@4:8I12c16", (superfunc)super_270, (IMP)meth_imp_270 },
	{ "@9@4:8^@12c16", (superfunc)super_271, (IMP)meth_imp_271 },
	{ "@9@4:8^v12c16", (superfunc)super_272, (IMP)meth_imp_272 },
	{ "@9@4:8^{OpaqueWindowPtr=}12c16", (superfunc)super_273, (IMP)meth_imp_273 },
	{ "@9@4:8^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}12c16", (superfunc)super_274, (IMP)meth_imp_274 },
	{ "@9@4:8^{_SelectionAnchor=iii}12c16", (superfunc)super_275, (IMP)meth_imp_275 },
	{ "@9@4:8c12c16", (superfunc)super_276, (IMP)meth_imp_276 },
	{ "@9@4:8i12c16", (superfunc)super_277, (IMP)meth_imp_277 },
	{ "C14@4:8I12^{OpaqueMenuHandle=}16S20", (superfunc)super_278, (IMP)meth_imp_278 },
	{ "C4@4:8", (superfunc)super_279, (IMP)meth_imp_279 },
	{ "I12@4:8:12@16", (superfunc)super_280, (IMP)meth_imp_280 },
	{ "I12@4:8@12@16", (superfunc)super_281, (IMP)meth_imp_281 },
	{ "I12@4:8@12I16", (superfunc)super_282, (IMP)meth_imp_282 },
	{ "I12@4:8I12*16", (superfunc)super_283, (IMP)meth_imp_283 },
	{ "I12@4:8I12^c16", (superfunc)super_284, (IMP)meth_imp_284 },
	{ "I12@4:8^I12@16", (superfunc)super_285, (IMP)meth_imp_285 },
	{ "I12@4:8r^v12I16", (superfunc)super_286, (IMP)meth_imp_286 },
	{ "I12@4:8{_NSPoint=ff}12", (superfunc)super_287, (IMP)meth_imp_287 },
	{ "I13@4:8@12@16c20", (superfunc)super_288, (IMP)meth_imp_288 },
	{ "I16@4:8@12@16@20", (superfunc)super_289, (IMP)meth_imp_289 },
	{ "I16@4:8@12{_NSRange=II}16", (superfunc)super_290, (IMP)meth_imp_290 },
	{ "I16@4:8^I12@16I20", (superfunc)super_291, (IMP)meth_imp_291 },
	{ "I16@4:8^I12{_NSRange=II}16", (superfunc)super_292, (IMP)meth_imp_292 },
	{ "I16@4:8{_NSPoint=ff}12@20", (superfunc)super_293, (IMP)meth_imp_293 },
	{ "I17@4:8@12i16@20c24", (superfunc)super_294, (IMP)meth_imp_294 },
	{ "I17@4:8@12{_NSRange=II}16c24", (superfunc)super_295, (IMP)meth_imp_295 },
	{ "I20@4:8^@12c16^@20@24", (superfunc)super_296, (IMP)meth_imp_296 },
	{ "I20@4:8{_NSPoint=ff}12@20^f24", (superfunc)super_297, (IMP)meth_imp_297 },
	{ "I24@4:8@12I16{_NSRange=II}20@28", (superfunc)super_298, (IMP)meth_imp_298 },
	{ "I28@4:8{_NSRange=II}12^I20^I24^i28^c32", (superfunc)super_299, (IMP)meth_imp_299 },
	{ "I4@4:8", (superfunc)super_300, (IMP)meth_imp_300 },
	{ "I5@4:8c12", (superfunc)super_301, (IMP)meth_imp_301 },
	{ "I6@4:8S12", (superfunc)super_302, (IMP)meth_imp_302 },
	{ "I8@4:8:12", (superfunc)super_303, (IMP)meth_imp_303 },
	{ "I8@4:8@12", (superfunc)super_304, (IMP)meth_imp_304 },
	{ "I8@4:8I12", (superfunc)super_305, (IMP)meth_imp_305 },
	{ "I8@4:8^I12", (superfunc)super_306, (IMP)meth_imp_306 },
	{ "I8@4:8^i12", (superfunc)super_307, (IMP)meth_imp_307 },
	{ "I8@4:8i12", (superfunc)super_308, (IMP)meth_imp_308 },
	{ "I8@4:8l12", (superfunc)super_309, (IMP)meth_imp_309 },
	{ "I9@4:8I12c16", (superfunc)super_310, (IMP)meth_imp_310 },
	{ "L4@4:8", (superfunc)super_311, (IMP)meth_imp_311 },
	{ "L8@4:8@12", (superfunc)super_312, (IMP)meth_imp_312 },
	{ "S4@4:8", (superfunc)super_313, (IMP)meth_imp_313 },
	{ "S8@4:8I12", (superfunc)super_314, (IMP)meth_imp_314 },
	{ "^*4@4:8", (superfunc)super_315, (IMP)meth_imp_315 },
	{ "^?8@4:8:12", (superfunc)super_316, (IMP)meth_imp_316 },
	{ "^S4@4:8", (superfunc)super_317, (IMP)meth_imp_317 },
	{ "^i12@4:8@12^i16", (superfunc)super_318, (IMP)meth_imp_318 },
	{ "^i4@4:8", (superfunc)super_319, (IMP)meth_imp_319 },
	{ "^i6@4:8S12", (superfunc)super_320, (IMP)meth_imp_320 },
	{ "^v12@4:8I12^{_NSRange=II}16", (superfunc)super_321, (IMP)meth_imp_321 },
	{ "^v20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12", (superfunc)super_322, (IMP)meth_imp_322 },
	{ "^v4@4:8", (superfunc)super_323, (IMP)meth_imp_323 },
	{ "^v5@4:8c12", (superfunc)super_324, (IMP)meth_imp_324 },
	{ "^v8@4:8@12", (superfunc)super_325, (IMP)meth_imp_325 },
	{ "^v8@4:8I12", (superfunc)super_326, (IMP)meth_imp_326 },
	{ "^v8@4:8^I12", (superfunc)super_327, (IMP)meth_imp_327 },
	{ "^{?=^{OpaquePMPrintSession}^{OpaquePMPrintSettings}^{OpaquePMPageFormat}}4@4:8", (superfunc)super_328, (IMP)meth_imp_328 },
	{ "^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12@4:8r*12^{?=b4b1b24(?=*^{?}^{__CFDictionary})}16", (superfunc)super_329, (IMP)meth_imp_329 },
	{ "^{?=b4b1b24(?=*^{?}^{__CFDictionary})}12@4:8r*12r*16", (superfunc)super_330, (IMP)meth_imp_330 },
	{ "^{?=b4b1b24(?=*^{?}^{__CFDictionary})}8@4:8i12", (superfunc)super_331, (IMP)meth_imp_331 },
	{ "^{AEDesc=I^^{OpaqueAEDataStorageType}}4@4:8", (superfunc)super_332, (IMP)meth_imp_332 },
	{ "^{CGFont=^{CGFontVTable}Ii^{CGEncoding}^{CGCMap}^{CGAdvanceSet}^{CGAdvanceSet}i^{CGFontCache}^vb1b1b1b1}4@4:8", (superfunc)super_333, (IMP)meth_imp_333 },
	{ "^{CGPDFDocument=}4@4:8", (superfunc)super_334, (IMP)meth_imp_334 },
	{ "^{ComponentInstanceRecord=[1l]}5@4:8c12", (superfunc)super_335, (IMP)meth_imp_335 },
	{ "^{FSRef=[80C]}4@4:8", (superfunc)super_336, (IMP)meth_imp_336 },
	{ "^{OpaqueCoreDragHandler=}4@4:8", (superfunc)super_337, (IMP)meth_imp_337 },
	{ "^{OpaqueGrafPtr=}4@4:8", (superfunc)super_338, (IMP)meth_imp_338 },
	{ "^{OpaqueIconRef=}4@4:8", (superfunc)super_339, (IMP)meth_imp_339 },
	{ "^{OpaquePMPageFormat=}4@4:8", (superfunc)super_340, (IMP)meth_imp_340 },
	{ "^{OpaquePMPrintSession=}4@4:8", (superfunc)super_341, (IMP)meth_imp_341 },
	{ "^{OpaquePMPrintSettings=}4@4:8", (superfunc)super_342, (IMP)meth_imp_342 },
	{ "^{OpaqueWindowPtr=}4@4:8", (superfunc)super_343, (IMP)meth_imp_343 },
	{ "^{_CoercerData=@:}12@4:8#12#16", (superfunc)super_344, (IMP)meth_imp_344 },
	{ "^{_NSFaceInfo=i^{_NSFaceInfo}@i{_NSFont_faceFlags=b1b1b1b1b1b1b1b1b1b1b22}^{_NSFontMetrics}^{_NSCGSFontMetrics}}8@4:8^{_NSFaceInfo=i^{_NSFaceInfo}@i{_NSFont_faceFlags=b1b1b1b1b1b1b1b1b1b1b22}^{_NSFontMetrics}^{_NSCGSFontMetrics}}12", (superfunc)super_345, (IMP)meth_imp_345 },
	{ "^{_NSMapTable=}5@4:8c12", (superfunc)super_346, (IMP)meth_imp_346 },
	{ "^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}12@4:8@12@16", (superfunc)super_347, (IMP)meth_imp_347 },
	{ "^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}24@4:8@12@16@20:24^v28", (superfunc)super_348, (IMP)meth_imp_348 },
	{ "^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}8@4:8@12", (superfunc)super_349, (IMP)meth_imp_349 },
	{ "^{_NSRect={_NSPoint=ff}{_NSSize=ff}}20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12", (superfunc)super_350, (IMP)meth_imp_350 },
	{ "^{_NSRect={_NSPoint=ff}{_NSSize=ff}}28@4:8{_NSRange=II}12{_NSRange=II}20@28^I32", (superfunc)super_351, (IMP)meth_imp_351 },
	{ "^{_NSRulebookSetHeader=i[4L]iiii[1i]}4@4:8", (superfunc)super_352, (IMP)meth_imp_352 },
	{ "^{_NSRulebookSetHeader=i[4L]iiii[1i]}8@4:8I12", (superfunc)super_353, (IMP)meth_imp_353 },
	{ "^{_NSRulebookTestStruct=iii[12i]}8@4:8I12", (superfunc)super_354, (IMP)meth_imp_354 },
	{ "^{_NSTypesetterGlyphInfo={_NSPoint=ff}fffI@{_NSSize=ff}{?=b1b1b1}}4@4:8", (superfunc)super_355, (IMP)meth_imp_355 },
	{ "^{_NSTypesetterGlyphInfo={_NSPoint=ff}fffI@{_NSSize=ff}{?=b1b1b1}}8@4:8i12", (superfunc)super_356, (IMP)meth_imp_356 },
	{ "^{_NSZone=}4@4:8", (superfunc)super_357, (IMP)meth_imp_357 },
	{ "^{_NXStream=I**iilii^{stream_functions}^v}4@4:8", (superfunc)super_358, (IMP)meth_imp_358 },
	{ "^{_PrivatePrintOperationInfo={_NSRect={_NSPoint=ff}{_NSSize=ff}}{_NSRect={_NSPoint=ff}{_NSSize=ff}}cccccccciiiiiii@@{_NSRect={_NSPoint=ff}{_NSSize=ff}}ccciffffii{_NSPoint=ff}I^{_NSModalSession}@iiciii@c@ic@@i@}4@4:8", (superfunc)super_359, (IMP)meth_imp_359 },
	{ "^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}12@4:8^{OpaqueIconRef=}12i16", (superfunc)super_360, (IMP)meth_imp_360 },
	{ "^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}16@4:8i12@16@20", (superfunc)super_361, (IMP)meth_imp_361 },
	{ "^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}32@4:8c12@16f36c24", (superfunc)super_362, (IMP)meth_imp_362 },
	{ "^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}8@4:8@12", (superfunc)super_363, (IMP)meth_imp_363 },
	{ "^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}12@4:8i12^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}16", (superfunc)super_364, (IMP)meth_imp_364 },
	{ "^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}13@4:8^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}12@16c20", (superfunc)super_365, (IMP)meth_imp_365 },
	{ "^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}20@4:8^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}12c16c20i24", (superfunc)super_366, (IMP)meth_imp_366 },
	{ "^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}8@4:8@12", (superfunc)super_367, (IMP)meth_imp_367 },
	{ "^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}8@4:8i12", (superfunc)super_368, (IMP)meth_imp_368 },
	{ "^{__CFArray=}5@4:8c12", (superfunc)super_369, (IMP)meth_imp_369 },
	{ "^{__CFArray=}8@4:8@12", (superfunc)super_370, (IMP)meth_imp_370 },
	{ "^{__CFDate=}4@4:8", (superfunc)super_371, (IMP)meth_imp_371 },
	{ "^{__CFDictionary=}8@4:8@12", (superfunc)super_372, (IMP)meth_imp_372 },
	{ "^{__CFHTTPMessage=}9@4:8@12c16", (superfunc)super_373, (IMP)meth_imp_373 },
	{ "^{__CFNotificationCenter=}4@4:8", (superfunc)super_374, (IMP)meth_imp_374 },
	{ "^{__CFPasteboard=}4@4:8", (superfunc)super_375, (IMP)meth_imp_375 },
	{ "^{__CFRunLoop=}4@4:8", (superfunc)super_376, (IMP)meth_imp_376 },
	{ "^{__CFSet=}5@4:8c12", (superfunc)super_377, (IMP)meth_imp_377 },
	{ "^{__CFSocket=}8@4:8@12", (superfunc)super_378, (IMP)meth_imp_378 },
	{ "^{__EventHandlerInfo=@:}12@4:8I12I16", (superfunc)super_379, (IMP)meth_imp_379 },
	{ "^{objc_method_description=:*}8@4:8:12", (superfunc)super_380, (IMP)meth_imp_380 },
	{ "c12@4:8#12@16", (superfunc)super_381, (IMP)meth_imp_381 },
	{ "c12@4:8*12I16", (superfunc)super_382, (IMP)meth_imp_382 },
	{ "c12@4:8:12@16", (superfunc)super_383, (IMP)meth_imp_383 },
	{ "c12@4:8@12:16", (superfunc)super_384, (IMP)meth_imp_384 },
	{ "c12@4:8@12@16", (superfunc)super_385, (IMP)meth_imp_385 },
	{ "c12@4:8@12I16", (superfunc)super_386, (IMP)meth_imp_386 },
	{ "c12@4:8@12^@16", (superfunc)super_387, (IMP)meth_imp_387 },
	{ "c12@4:8@12^c16", (superfunc)super_388, (IMP)meth_imp_388 },
	{ "c12@4:8@12^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}16", (superfunc)super_389, (IMP)meth_imp_389 },
	{ "c12@4:8@12i16", (superfunc)super_390, (IMP)meth_imp_390 },
	{ "c12@4:8@12r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_391, (IMP)meth_imp_391 },
	{ "c12@4:8I12I16", (superfunc)super_392, (IMP)meth_imp_392 },
	{ "c12@4:8^@12@16", (superfunc)super_393, (IMP)meth_imp_393 },
	{ "c12@4:8^@12I16", (superfunc)super_394, (IMP)meth_imp_394 },
	{ "c12@4:8^@12^I16", (superfunc)super_395, (IMP)meth_imp_395 },
	{ "c12@4:8^{FSRef=[80C]}12@16", (superfunc)super_396, (IMP)meth_imp_396 },
	{ "c12@4:8^{tiff=*^{_NXStream}sccsll{?=IIIIIISSSSSSSSSSIIIffSSffII[2S]ISSSSI^S^S^S^S[3^S]*********[2I]II^I^I[2S]^f[2S]S^f^f^f[4^S]S[2S]**I^v}{?=SSL}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}12i16", (superfunc)super_397, (IMP)meth_imp_397 },
	{ "c12@4:8i12@16", (superfunc)super_398, (IMP)meth_imp_398 },
	{ "c12@4:8i12i16", (superfunc)super_399, (IMP)meth_imp_399 },
	{ "c12@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@16", (superfunc)super_400, (IMP)meth_imp_400 },
	{ "c12@4:8{NSButtonState=iccc}12", (superfunc)super_401, (IMP)meth_imp_401 },
	{ "c12@4:8{_NSPoint=ff}12", (superfunc)super_402, (IMP)meth_imp_402 },
	{ "c13@4:8@12@16c20", (superfunc)super_403, (IMP)meth_imp_403 },
	{ "c13@4:8@12c16c20", (superfunc)super_404, (IMP)meth_imp_404 },
	{ "c14@4:8@12@16S20", (superfunc)super_405, (IMP)meth_imp_405 },
	{ "c16@4:8*12I16@20", (superfunc)super_406, (IMP)meth_imp_406 },
	{ "c16@4:8*12I16I20", (superfunc)super_407, (IMP)meth_imp_407 },
	{ "c16@4:8:12@16@20", (superfunc)super_408, (IMP)meth_imp_408 },
	{ "c16@4:8@12@16:20", (superfunc)super_409, (IMP)meth_imp_409 },
	{ "c16@4:8@12@16@20", (superfunc)super_410, (IMP)meth_imp_410 },
	{ "c16@4:8@12@16I20", (superfunc)super_411, (IMP)meth_imp_411 },
	{ "c16@4:8@12@16^c20", (superfunc)super_412, (IMP)meth_imp_412 },
	{ "c16@4:8@12@16i20", (superfunc)super_413, (IMP)meth_imp_413 },
	{ "c16@4:8@12^@16^@20", (superfunc)super_414, (IMP)meth_imp_414 },
	{ "c16@4:8@12^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16^c20", (superfunc)super_415, (IMP)meth_imp_415 },
	{ "c16@4:8@12i16i20", (superfunc)super_416, (IMP)meth_imp_416 },
	{ "c16@4:8@12r^{FSRef=[80C]}16r^{FSRef=[80C]}20", (superfunc)super_417, (IMP)meth_imp_417 },
	{ "c16@4:8@12r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16i20", (superfunc)super_418, (IMP)meth_imp_418 },
	{ "c16@4:8@12{_NSPoint=ff}16", (superfunc)super_419, (IMP)meth_imp_419 },
	{ "c16@4:8@12{_NSRange=II}16", (superfunc)super_420, (IMP)meth_imp_420 },
	{ "c16@4:8I12I16@20", (superfunc)super_421, (IMP)meth_imp_421 },
	{ "c16@4:8^@12@16^@20", (superfunc)super_422, (IMP)meth_imp_422 },
	{ "c16@4:8^I12^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@20", (superfunc)super_423, (IMP)meth_imp_423 },
	{ "c16@4:8^i12^i16@20", (superfunc)super_424, (IMP)meth_imp_424 },
	{ "c16@4:8i12@16@20", (superfunc)super_425, (IMP)meth_imp_425 },
	{ "c16@4:8i12i16i20", (superfunc)super_426, (IMP)meth_imp_426 },
	{ "c16@4:8s12r^{FSRef=[80C]}16^{FSRef=[80C]}20", (superfunc)super_427, (IMP)meth_imp_427 },
	{ "c16@4:8{_NSPoint=ff}12@20", (superfunc)super_428, (IMP)meth_imp_428 },
	{ "c16@4:8{_NSPoint=ff}12i20", (superfunc)super_429, (IMP)meth_imp_429 },
	{ "c17@4:8@12^{FSRef=[80C]}16c20c24", (superfunc)super_430, (IMP)meth_imp_430 },
	{ "c20@4:8:12@16i20i24", (superfunc)super_431, (IMP)meth_imp_431 },
	{ "c20@4:8@12@16@20I24", (superfunc)super_432, (IMP)meth_imp_432 },
	{ "c20@4:8@12@16@20i24", (superfunc)super_433, (IMP)meth_imp_433 },
	{ "c20@4:8@12{_NSRange=II}16@24", (superfunc)super_434, (IMP)meth_imp_434 },
	{ "c20@4:8^@12@16I20@24", (superfunc)super_435, (IMP)meth_imp_435 },
	{ "c20@4:8^i12^i16@20r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}24", (superfunc)super_436, (IMP)meth_imp_436 },
	{ "c20@4:8^i12^i16{_NSPoint=ff}20", (superfunc)super_437, (IMP)meth_imp_437 },
	{ "c20@4:8i12@16@20@24", (superfunc)super_438, (IMP)meth_imp_438 },
	{ "c20@4:8{_NSPoint=ff}12^i20^i24", (superfunc)super_439, (IMP)meth_imp_439 },
	{ "c20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12", (superfunc)super_440, (IMP)meth_imp_440 },
	{ "c21@4:8*12i16c20c24c28", (superfunc)super_441, (IMP)meth_imp_441 },
	{ "c21@4:8@12@16c20c24c28", (superfunc)super_442, (IMP)meth_imp_442 },
	{ "c21@4:8@12I16^@20@24c28", (superfunc)super_443, (IMP)meth_imp_443 },
	{ "c24@4:8@12@16@20@24^i28", (superfunc)super_444, (IMP)meth_imp_444 },
	{ "c24@4:8@12@16i20^{_NSMapTable=}24@28", (superfunc)super_445, (IMP)meth_imp_445 },
	{ "c24@4:8@12@16{_NSPoint=ff}20@28", (superfunc)super_446, (IMP)meth_imp_446 },
	{ "c24@4:8@12I16@20@24I28", (superfunc)super_447, (IMP)meth_imp_447 },
	{ "c24@4:8@12i16^c20^c24^@28", (superfunc)super_448, (IMP)meth_imp_448 },
	{ "c24@4:8@12r^{FSRef=[80C]}16r^{FSRef=[80C]}20@24i28", (superfunc)super_449, (IMP)meth_imp_449 },
	{ "c24@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_450, (IMP)meth_imp_450 },
	{ "c24@4:8I12{_NSPoint=ff}16I24@28", (superfunc)super_451, (IMP)meth_imp_451 },
	{ "c24@4:8{_NSPoint=ff}12{_NSPoint=ff}20@28", (superfunc)super_452, (IMP)meth_imp_452 },
	{ "c24@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28", (superfunc)super_453, (IMP)meth_imp_453 },
	{ "c25@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16c32", (superfunc)super_454, (IMP)meth_imp_454 },
	{ "c25@4:8^i12@16@20i24c28c32", (superfunc)super_455, (IMP)meth_imp_455 },
	{ "c28@4:8@12^c16^c20^c24^@28^@32", (superfunc)super_456, (IMP)meth_imp_456 },
	{ "c28@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32", (superfunc)super_457, (IMP)meth_imp_457 },
	{ "c28@4:8^@12^{_NSRange=II}16@20{_NSRange=II}24^@32", (superfunc)super_458, (IMP)meth_imp_458 },
	{ "c28@4:8{_NSPoint=ff}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}20", (superfunc)super_459, (IMP)meth_imp_459 },
	{ "c28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32", (superfunc)super_460, (IMP)meth_imp_460 },
	{ "c32@4:8^i12{_NSSize=ff}16f36", (superfunc)super_461, (IMP)meth_imp_461 },
	{ "c32@4:8f36", (superfunc)super_462, (IMP)meth_imp_462 },
	{ "c32@4:8f36c16", (superfunc)super_463, (IMP)meth_imp_463 },
	{ "c32@4:8i12f36r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}20r^{_NSPoint=ff}24", (superfunc)super_464, (IMP)meth_imp_464 },
	{ "c32@4:8r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12f36", (superfunc)super_465, (IMP)meth_imp_465 },
	{ "c36@4:8@12^{FSRef=[80C]}16@20^{FSRef=[80C]}24i28^{_NSMapTable=}32@40", (superfunc)super_466, (IMP)meth_imp_466 },
	{ "c36@4:8@12i16i20c24c28c32c43", (superfunc)super_467, (IMP)meth_imp_467 },
	{ "c36@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32I40", (superfunc)super_468, (IMP)meth_imp_468 },
	{ "c36@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32c43", (superfunc)super_469, (IMP)meth_imp_469 },
	{ "c36@4:8d36", (superfunc)super_470, (IMP)meth_imp_470 },
	{ "c36@4:8d36^v20@24@28I32", (superfunc)super_471, (IMP)meth_imp_471 },
	{ "c36@4:8{_NSRange=II}12{_NSRange=II}20{_NSRange=II}28@40", (superfunc)super_472, (IMP)meth_imp_472 },
	{ "c36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28i32i40", (superfunc)super_473, (IMP)meth_imp_473 },
	{ "c40@4:8*12I16^I20I24c28{_NSRange=II}36^{_NSRange=II}44", (superfunc)super_474, (IMP)meth_imp_474 },
	{ "c40@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32I40c47", (superfunc)super_475, (IMP)meth_imp_475 },
	{ "c40@4:8^@12I16^I20I24c28{_NSRange=II}36^{_NSRange=II}44", (superfunc)super_476, (IMP)meth_imp_476 },
	{ "c40@4:8d36@20@24@28@32I40I44", (superfunc)super_477, (IMP)meth_imp_477 },
	{ "c4@4:8", (superfunc)super_478, (IMP)meth_imp_478 },
	{ "c56@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32i48f36c59c63", (superfunc)super_479, (IMP)meth_imp_479 },
	{ "c5@4:8c12", (superfunc)super_480, (IMP)meth_imp_480 },
	{ "c6@4:8S12", (superfunc)super_481, (IMP)meth_imp_481 },
	{ "c6@4:8s12", (superfunc)super_482, (IMP)meth_imp_482 },
	{ "c8@4:8#12", (superfunc)super_483, (IMP)meth_imp_483 },
	{ "c8@4:8:12", (superfunc)super_484, (IMP)meth_imp_484 },
	{ "c8@4:8@12", (superfunc)super_485, (IMP)meth_imp_485 },
	{ "c8@4:8I12", (superfunc)super_486, (IMP)meth_imp_486 },
	{ "c8@4:8L12", (superfunc)super_487, (IMP)meth_imp_487 },
	{ "c8@4:8^*12", (superfunc)super_488, (IMP)meth_imp_488 },
	{ "c8@4:8^I12", (superfunc)super_489, (IMP)meth_imp_489 },
	{ "c8@4:8^d12", (superfunc)super_490, (IMP)meth_imp_490 },
	{ "c8@4:8^f12", (superfunc)super_491, (IMP)meth_imp_491 },
	{ "c8@4:8^i12", (superfunc)super_492, (IMP)meth_imp_492 },
	{ "c8@4:8^q12", (superfunc)super_493, (IMP)meth_imp_493 },
	{ "c8@4:8^v12", (superfunc)super_494, (IMP)meth_imp_494 },
	{ "c8@4:8^{_NSPoint=ff}12", (superfunc)super_495, (IMP)meth_imp_495 },
	{ "c8@4:8^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}12", (superfunc)super_496, (IMP)meth_imp_496 },
	{ "c8@4:8i12", (superfunc)super_497, (IMP)meth_imp_497 },
	{ "c8@4:8r*12", (superfunc)super_498, (IMP)meth_imp_498 },
	{ "c8@4:8r^{FSRef=[80C]}12", (superfunc)super_499, (IMP)meth_imp_499 },
	{ "c8@4:8r^{_NSPoint=ff}12", (superfunc)super_500, (IMP)meth_imp_500 },
	{ "c9@4:8@12c16", (superfunc)super_501, (IMP)meth_imp_501 },
	{ "c9@4:8^{_NSPoint=ff}12c16", (superfunc)super_502, (IMP)meth_imp_502 },
	{ "c9@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c16", (superfunc)super_503, (IMP)meth_imp_503 },
	{ "c9@4:8^{_NSSize=ff}12c16", (superfunc)super_504, (IMP)meth_imp_504 },
	{ "c9@4:8^{_RepresentationInfo=^{_RepresentationInfo}^{_CacheWindowInfo}{_CacheRect=SSSS}@{_RepresentationInfoFlags=b1b1b1b4b1b24}@@^vi}12c16", (superfunc)super_505, (IMP)meth_imp_505 },
	{ "c9@4:8i12c16", (superfunc)super_506, (IMP)meth_imp_506 },
	{ "d20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12", (superfunc)super_507, (IMP)meth_imp_507 },
	{ "d36@4:8d36", (superfunc)super_508, (IMP)meth_imp_508 },
	{ "d4@4:8", (superfunc)super_509, (IMP)meth_imp_509 },
	{ "d8@4:8@12", (superfunc)super_510, (IMP)meth_imp_510 },
	{ "d8@4:8i12", (superfunc)super_511, (IMP)meth_imp_511 },
	{ "f12@4:8@12@16", (superfunc)super_512, (IMP)meth_imp_512 },
	{ "f12@4:8@12I16", (superfunc)super_513, (IMP)meth_imp_513 },
	{ "f12@4:8r*12I16", (superfunc)super_514, (IMP)meth_imp_514 },
	{ "f12@4:8{_NSSize=ff}12", (superfunc)super_515, (IMP)meth_imp_515 },
	{ "f16@4:8{_NSPoint=ff}12@20", (superfunc)super_516, (IMP)meth_imp_516 },
	{ "f32@4:8@12@16f36", (superfunc)super_517, (IMP)meth_imp_517 },
	{ "f32@4:8c12f36", (superfunc)super_518, (IMP)meth_imp_518 },
	{ "f32@4:8f36", (superfunc)super_519, (IMP)meth_imp_519 },
	{ "f36@4:8d36", (superfunc)super_520, (IMP)meth_imp_520 },
	{ "f4@4:8", (superfunc)super_521, (IMP)meth_imp_521 },
	{ "f8@4:8@12", (superfunc)super_522, (IMP)meth_imp_522 },
	{ "f8@4:8I12", (superfunc)super_523, (IMP)meth_imp_523 },
	{ "f8@4:8i12", (superfunc)super_524, (IMP)meth_imp_524 },
	{ "i12@4:8*12@16", (superfunc)super_525, (IMP)meth_imp_525 },
	{ "i12@4:8@12:16", (superfunc)super_526, (IMP)meth_imp_526 },
	{ "i12@4:8@12@16", (superfunc)super_527, (IMP)meth_imp_527 },
	{ "i12@4:8@12I16", (superfunc)super_528, (IMP)meth_imp_528 },
	{ "i12@4:8@12^i16", (superfunc)super_529, (IMP)meth_imp_529 },
	{ "i12@4:8@12i16", (superfunc)super_530, (IMP)meth_imp_530 },
	{ "i12@4:8S12i16", (superfunc)super_531, (IMP)meth_imp_531 },
	{ "i12@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12^f16", (superfunc)super_532, (IMP)meth_imp_532 },
	{ "i12@4:8^{__sFILE=*iiss{__sbuf=*i}i^v^?^?^?^?{__sbuf=*i}*i[3C][1C]{__sbuf=*i}iq}12i16", (superfunc)super_533, (IMP)meth_imp_533 },
	{ "i12@4:8i12@16", (superfunc)super_534, (IMP)meth_imp_534 },
	{ "i12@4:8i12I16", (superfunc)super_535, (IMP)meth_imp_535 },
	{ "i12@4:8i12^{_NSPoint=ff}16", (superfunc)super_536, (IMP)meth_imp_536 },
	{ "i12@4:8i12i16", (superfunc)super_537, (IMP)meth_imp_537 },
	{ "i12@4:8r*12^i16", (superfunc)super_538, (IMP)meth_imp_538 },
	{ "i12@4:8{NSButtonState=iccc}12", (superfunc)super_539, (IMP)meth_imp_539 },
	{ "i12@4:8{_NSPoint=ff}12", (superfunc)super_540, (IMP)meth_imp_540 },
	{ "i13@4:8@12@16c20", (superfunc)super_541, (IMP)meth_imp_541 },
	{ "i13@4:8@12i16c20", (superfunc)super_542, (IMP)meth_imp_542 },
	{ "i16@4:8@12@16@20", (superfunc)super_543, (IMP)meth_imp_543 },
	{ "i16@4:8@12@16i20", (superfunc)super_544, (IMP)meth_imp_544 },
	{ "i16@4:8@12c16@20", (superfunc)super_545, (IMP)meth_imp_545 },
	{ "i16@4:8@12{_NSRange=II}16", (superfunc)super_546, (IMP)meth_imp_546 },
	{ "i16@4:8^I12i16^{_NSPoint=ff}20", (superfunc)super_547, (IMP)meth_imp_547 },
	{ "i16@4:8i12c16@20", (superfunc)super_548, (IMP)meth_imp_548 },
	{ "i16@4:8i12i16@20", (superfunc)super_549, (IMP)meth_imp_549 },
	{ "i16@4:8i12{_NSPoint=ff}16", (superfunc)super_550, (IMP)meth_imp_550 },
	{ "i17@4:8@12@16@20c24", (superfunc)super_551, (IMP)meth_imp_551 },
	{ "i20@4:8@12@16@20@24", (superfunc)super_552, (IMP)meth_imp_552 },
	{ "i20@4:8@12I16{_NSRange=II}20", (superfunc)super_553, (IMP)meth_imp_553 },
	{ "i20@4:8@12^S16^i20^{_NSSortState=iIIII[4@]}24", (superfunc)super_554, (IMP)meth_imp_554 },
	{ "i20@4:8^{OpaqueEventRef=}12{Point=ss}16s20I24", (superfunc)super_555, (IMP)meth_imp_555 },
	{ "i20@4:8c12@16@20@24", (superfunc)super_556, (IMP)meth_imp_556 },
	{ "i20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12", (superfunc)super_557, (IMP)meth_imp_557 },
	{ "i24@4:8@12@16@20@24^@28", (superfunc)super_558, (IMP)meth_imp_558 },
	{ "i24@4:8@12I16{_NSRange=II}20@28", (superfunc)super_559, (IMP)meth_imp_559 },
	{ "i24@4:8@12c16@20@24@28", (superfunc)super_560, (IMP)meth_imp_560 },
	{ "i24@4:8i12{_NSPoint=ff}16@24i28", (superfunc)super_561, (IMP)meth_imp_561 },
	{ "i28@4:8@12@16@20@24@28@32", (superfunc)super_562, (IMP)meth_imp_562 },
	{ "i28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28^v32", (superfunc)super_563, (IMP)meth_imp_563 },
	{ "i32@4:8f36", (superfunc)super_564, (IMP)meth_imp_564 },
	{ "i32@4:8i12f36", (superfunc)super_565, (IMP)meth_imp_565 },
	{ "i36@4:8@12@16i20c24c28c32c43", (superfunc)super_566, (IMP)meth_imp_566 },
	{ "i36@4:8@12{_NSRange=II}16@24{_NSRange=II}28i40", (superfunc)super_567, (IMP)meth_imp_567 },
	{ "i36@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32^v40", (superfunc)super_568, (IMP)meth_imp_568 },
	{ "i36@4:8d36", (superfunc)super_569, (IMP)meth_imp_569 },
	{ "i36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28^v32c43", (superfunc)super_570, (IMP)meth_imp_570 },
	{ "i36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28@32^v40", (superfunc)super_571, (IMP)meth_imp_571 },
	{ "i40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28@32@40@44", (superfunc)super_572, (IMP)meth_imp_572 },
	{ "i48@4:8@12@16@20{_NSRect={_NSPoint=ff}{_NSSize=ff}}28@44c51^v52", (superfunc)super_573, (IMP)meth_imp_573 },
	{ "i4@4:8", (superfunc)super_574, (IMP)meth_imp_574 },
	{ "i5@4:8c12", (superfunc)super_575, (IMP)meth_imp_575 },
	{ "i6@4:8S12", (superfunc)super_576, (IMP)meth_imp_576 },
	{ "i8@4:8*12", (superfunc)super_577, (IMP)meth_imp_577 },
	{ "i8@4:8@12", (superfunc)super_578, (IMP)meth_imp_578 },
	{ "i8@4:8I12", (superfunc)super_579, (IMP)meth_imp_579 },
	{ "i8@4:8^@12", (superfunc)super_580, (IMP)meth_imp_580 },
	{ "i8@4:8^I12", (superfunc)super_581, (IMP)meth_imp_581 },
	{ "i8@4:8^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}12", (superfunc)super_582, (IMP)meth_imp_582 },
	{ "i8@4:8i12", (superfunc)super_583, (IMP)meth_imp_583 },
	{ "i8@4:8r^{_NSPoint=ff}12", (superfunc)super_584, (IMP)meth_imp_584 },
	{ "i9@4:8@12c16", (superfunc)super_585, (IMP)meth_imp_585 },
	{ "l4@4:8", (superfunc)super_586, (IMP)meth_imp_586 },
	{ "q4@4:8", (superfunc)super_587, (IMP)meth_imp_587 },
	{ "q8@4:8@12", (superfunc)super_588, (IMP)meth_imp_588 },
	{ "r*4@4:8", (superfunc)super_589, (IMP)meth_imp_589 },
	{ "r*5@4:8c12", (superfunc)super_590, (IMP)meth_imp_590 },
	{ "r*8@4:8@12", (superfunc)super_591, (IMP)meth_imp_591 },
	{ "r*8@4:8I12", (superfunc)super_592, (IMP)meth_imp_592 },
	{ "r^I4@4:8", (superfunc)super_593, (IMP)meth_imp_593 },
	{ "r^f4@4:8", (superfunc)super_594, (IMP)meth_imp_594 },
	{ "r^f8@4:8@12", (superfunc)super_595, (IMP)meth_imp_595 },
	{ "r^i4@4:8", (superfunc)super_596, (IMP)meth_imp_596 },
	{ "r^v4@4:8", (superfunc)super_597, (IMP)meth_imp_597 },
	{ "r^{FSRef=[80C]}4@4:8", (superfunc)super_598, (IMP)meth_imp_598 },
	{ "s12@4:8@12@16", (superfunc)super_599, (IMP)meth_imp_599 },
	{ "s12@4:8L12@16", (superfunc)super_600, (IMP)meth_imp_600 },
	{ "s16@4:8@12@16@20", (superfunc)super_601, (IMP)meth_imp_601 },
	{ "s16@4:8L12@16@20", (superfunc)super_602, (IMP)meth_imp_602 },
	{ "s16@4:8r^{AEDesc=I^^{OpaqueAEDataStorageType}}12^{AEDesc=I^^{OpaqueAEDataStorageType}}16I20", (superfunc)super_603, (IMP)meth_imp_603 },
	{ "s4@4:8", (superfunc)super_604, (IMP)meth_imp_604 },
	{ "s8@4:8@12", (superfunc)super_605, (IMP)meth_imp_605 },
	{ "v104@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32{_NSRect={_NSPoint=ff}{_NSSize=ff}}48{_NSRect={_NSPoint=ff}{_NSSize=ff}}64{_NSRect={_NSPoint=ff}{_NSSize=ff}}80{_NSRect={_NSPoint=ff}{_NSSize=ff}}96", (superfunc)super_606, (IMP)meth_imp_606 },
	{ "v10@4:8@12s16", (superfunc)super_607, (IMP)meth_imp_607 },
	{ "v10@4:8^{OpaqueIconRef=}12s16", (superfunc)super_608, (IMP)meth_imp_608 },
	{ "v12@4:8#12^v16", (superfunc)super_609, (IMP)meth_imp_609 },
	{ "v12@4:8*12I16", (superfunc)super_610, (IMP)meth_imp_610 },
	{ "v12@4:8:12@16", (superfunc)super_611, (IMP)meth_imp_611 },
	{ "v12@4:8@12#16", (superfunc)super_612, (IMP)meth_imp_612 },
	{ "v12@4:8@12:16", (superfunc)super_613, (IMP)meth_imp_613 },
	{ "v12@4:8@12@16", (superfunc)super_614, (IMP)meth_imp_614 },
	{ "v12@4:8@12I16", (superfunc)super_615, (IMP)meth_imp_615 },
	{ "v12@4:8@12L16", (superfunc)super_616, (IMP)meth_imp_616 },
	{ "v12@4:8@12^c16", (superfunc)super_617, (IMP)meth_imp_617 },
	{ "v12@4:8@12^i16", (superfunc)super_618, (IMP)meth_imp_618 },
	{ "v12@4:8@12^v16", (superfunc)super_619, (IMP)meth_imp_619 },
	{ "v12@4:8@12^{?=^SI^SI^SI}16", (superfunc)super_620, (IMP)meth_imp_620 },
	{ "v12@4:8@12i16", (superfunc)super_621, (IMP)meth_imp_621 },
	{ "v12@4:8@12l16", (superfunc)super_622, (IMP)meth_imp_622 },
	{ "v12@4:8@16", (superfunc)super_623, (IMP)meth_imp_623 },
	{ "v12@4:8I12@16", (superfunc)super_624, (IMP)meth_imp_624 },
	{ "v12@4:8I12I16", (superfunc)super_625, (IMP)meth_imp_625 },
	{ "v12@4:8I12^v16", (superfunc)super_626, (IMP)meth_imp_626 },
	{ "v12@4:8Q12", (superfunc)super_627, (IMP)meth_imp_627 },
	{ "v12@4:8S12I16", (superfunc)super_628, (IMP)meth_imp_628 },
	{ "v12@4:8^?12^v16", (superfunc)super_629, (IMP)meth_imp_629 },
	{ "v12@4:8^@12^@16", (superfunc)super_630, (IMP)meth_imp_630 },
	{ "v12@4:8^@12^i16", (superfunc)super_631, (IMP)meth_imp_631 },
	{ "v12@4:8^@12^{_NSRange=II}16", (superfunc)super_632, (IMP)meth_imp_632 },
	{ "v12@4:8^@12^{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_633, (IMP)meth_imp_633 },
	{ "v12@4:8^I12I16", (superfunc)super_634, (IMP)meth_imp_634 },
	{ "v12@4:8^I12^I16", (superfunc)super_635, (IMP)meth_imp_635 },
	{ "v12@4:8^^S12^i16", (superfunc)super_636, (IMP)meth_imp_636 },
	{ "v12@4:8^^{OpaqueIconRef}12^s16", (superfunc)super_637, (IMP)meth_imp_637 },
	{ "v12@4:8^f12^f16", (superfunc)super_638, (IMP)meth_imp_638 },
	{ "v12@4:8^i12I16", (superfunc)super_639, (IMP)meth_imp_639 },
	{ "v12@4:8^i12^f16", (superfunc)super_640, (IMP)meth_imp_640 },
	{ "v12@4:8^i12^i16", (superfunc)super_641, (IMP)meth_imp_641 },
	{ "v12@4:8^l12i16", (superfunc)super_642, (IMP)meth_imp_642 },
	{ "v12@4:8^v12I16", (superfunc)super_643, (IMP)meth_imp_643 },
	{ "v12@4:8^v12i16", (superfunc)super_644, (IMP)meth_imp_644 },
	{ "v12@4:8^{_NSPoint=ff}12i16", (superfunc)super_645, (IMP)meth_imp_645 },
	{ "v12@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12i16", (superfunc)super_646, (IMP)meth_imp_646 },
	{ "v12@4:8^{_RowEntry=^{_RowEntry}^{_RowEntry}@sscccc}12i16", (superfunc)super_647, (IMP)meth_imp_647 },
	{ "v12@4:8^{__CFReadStream=}12@16", (superfunc)super_648, (IMP)meth_imp_648 },
	{ "v12@4:8c12@16", (superfunc)super_649, (IMP)meth_imp_649 },
	{ "v12@4:8c12I16", (superfunc)super_650, (IMP)meth_imp_650 },
	{ "v12@4:8i12@16", (superfunc)super_651, (IMP)meth_imp_651 },
	{ "v12@4:8i12I16", (superfunc)super_652, (IMP)meth_imp_652 },
	{ "v12@4:8i12i16", (superfunc)super_653, (IMP)meth_imp_653 },
	{ "v12@4:8r*12^v16", (superfunc)super_654, (IMP)meth_imp_654 },
	{ "v12@4:8r*12i16", (superfunc)super_655, (IMP)meth_imp_655 },
	{ "v12@4:8r*12r^v16", (superfunc)super_656, (IMP)meth_imp_656 },
	{ "v12@4:8r*16", (superfunc)super_657, (IMP)meth_imp_657 },
	{ "v12@4:8r^S12i16", (superfunc)super_658, (IMP)meth_imp_658 },
	{ "v12@4:8r^^i12^i16", (superfunc)super_659, (IMP)meth_imp_659 },
	{ "v12@4:8r^i12i16", (superfunc)super_660, (IMP)meth_imp_660 },
	{ "v12@4:8r^v12I16", (superfunc)super_661, (IMP)meth_imp_661 },
	{ "v12@4:8r^{_NSPoint=ff}12@16", (superfunc)super_662, (IMP)meth_imp_662 },
	{ "v12@4:8{_NSPoint=ff}12", (superfunc)super_663, (IMP)meth_imp_663 },
	{ "v12@4:8{_NSRange=II}12", (superfunc)super_664, (IMP)meth_imp_664 },
	{ "v12@4:8{_NSSize=ff}12", (superfunc)super_665, (IMP)meth_imp_665 },
	{ "v13@4:8:12@16c20", (superfunc)super_666, (IMP)meth_imp_666 },
	{ "v13@4:8@12@16c20", (superfunc)super_667, (IMP)meth_imp_667 },
	{ "v13@4:8@12^i16c20", (superfunc)super_668, (IMP)meth_imp_668 },
	{ "v13@4:8@12c16c20", (superfunc)super_669, (IMP)meth_imp_669 },
	{ "v13@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@16c20", (superfunc)super_670, (IMP)meth_imp_670 },
	{ "v13@4:8i12c16c20", (superfunc)super_671, (IMP)meth_imp_671 },
	{ "v13@4:8i12i16c20", (superfunc)super_672, (IMP)meth_imp_672 },
	{ "v13@4:8{_NSRange=II}12c20", (superfunc)super_673, (IMP)meth_imp_673 },
	{ "v16@4:8:12@16@20", (superfunc)super_674, (IMP)meth_imp_674 },
	{ "v16@4:8:12i16i20", (superfunc)super_675, (IMP)meth_imp_675 },
	{ "v16@4:8@12:16#20", (superfunc)super_676, (IMP)meth_imp_676 },
	{ "v16@4:8@12:16@20", (superfunc)super_677, (IMP)meth_imp_677 },
	{ "v16@4:8@12:16I20", (superfunc)super_678, (IMP)meth_imp_678 },
	{ "v16@4:8@12:16^v20", (superfunc)super_679, (IMP)meth_imp_679 },
	{ "v16@4:8@12@16*20", (superfunc)super_680, (IMP)meth_imp_680 },
	{ "v16@4:8@12@16@20", (superfunc)super_681, (IMP)meth_imp_681 },
	{ "v16@4:8@12@16I20", (superfunc)super_682, (IMP)meth_imp_682 },
	{ "v16@4:8@12@16L20", (superfunc)super_683, (IMP)meth_imp_683 },
	{ "v16@4:8@12@16i20", (superfunc)super_684, (IMP)meth_imp_684 },
	{ "v16@4:8@12@20", (superfunc)super_685, (IMP)meth_imp_685 },
	{ "v16@4:8@12I16@20", (superfunc)super_686, (IMP)meth_imp_686 },
	{ "v16@4:8@12^@16^@20", (superfunc)super_687, (IMP)meth_imp_687 },
	{ "v16@4:8@12c16^v20", (superfunc)super_688, (IMP)meth_imp_688 },
	{ "v16@4:8@12i16@20", (superfunc)super_689, (IMP)meth_imp_689 },
	{ "v16@4:8@12i16I20", (superfunc)super_690, (IMP)meth_imp_690 },
	{ "v16@4:8@12i16^v20", (superfunc)super_691, (IMP)meth_imp_691 },
	{ "v16@4:8@12i16i20", (superfunc)super_692, (IMP)meth_imp_692 },
	{ "v16@4:8@12{_NSPoint=ff}16", (superfunc)super_693, (IMP)meth_imp_693 },
	{ "v16@4:8@12{_NSRange=II}16", (superfunc)super_694, (IMP)meth_imp_694 },
	{ "v16@4:8@12{_NSSize=ff}16", (superfunc)super_695, (IMP)meth_imp_695 },
	{ "v16@4:8I12@16@20", (superfunc)super_696, (IMP)meth_imp_696 },
	{ "v16@4:8I12I16I20", (superfunc)super_697, (IMP)meth_imp_697 },
	{ "v16@4:8I12^v16L20", (superfunc)super_698, (IMP)meth_imp_698 },
	{ "v16@4:8^@12{_NSRange=II}16", (superfunc)super_699, (IMP)meth_imp_699 },
	{ "v16@4:8^I12i16@20", (superfunc)super_700, (IMP)meth_imp_700 },
	{ "v16@4:8^S12^i16^{?=^SI^SI^SI}20", (superfunc)super_701, (IMP)meth_imp_701 },
	{ "v16@4:8^S12{_NSRange=II}16", (superfunc)super_702, (IMP)meth_imp_702 },
	{ "v16@4:8^^{OpaqueIconRef}12^s16@20", (superfunc)super_703, (IMP)meth_imp_703 },
	{ "v16@4:8^f12^i16^f20", (superfunc)super_704, (IMP)meth_imp_704 },
	{ "v16@4:8^i12I16I20", (superfunc)super_705, (IMP)meth_imp_705 },
	{ "v16@4:8^i12I16^I20", (superfunc)super_706, (IMP)meth_imp_706 },
	{ "v16@4:8^l12i16i20", (superfunc)super_707, (IMP)meth_imp_707 },
	{ "v16@4:8^v12I16I20", (superfunc)super_708, (IMP)meth_imp_708 },
	{ "v16@4:8^v12I16^I20", (superfunc)super_709, (IMP)meth_imp_709 },
	{ "v16@4:8^v12{_NSRange=II}16", (superfunc)super_710, (IMP)meth_imp_710 },
	{ "v16@4:8^{_NSMapTable=}12r*16@20", (superfunc)super_711, (IMP)meth_imp_711 },
	{ "v16@4:8^{__CFData=}12^{__CFData=}16^{__CFSocket=}20", (superfunc)super_712, (IMP)meth_imp_712 },
	{ "v16@4:8^{__CFString=}12I16I20", (superfunc)super_713, (IMP)meth_imp_713 },
	{ "v16@4:8c12I16I20", (superfunc)super_714, (IMP)meth_imp_714 },
	{ "v16@4:8c12i16i20", (superfunc)super_715, (IMP)meth_imp_715 },
	{ "v16@4:8c12{_NSPoint=ff}16", (superfunc)super_716, (IMP)meth_imp_716 },
	{ "v16@4:8i12Q16", (superfunc)super_717, (IMP)meth_imp_717 },
	{ "v16@4:8i12i16@20", (superfunc)super_718, (IMP)meth_imp_718 },
	{ "v16@4:8i12i16I20", (superfunc)super_719, (IMP)meth_imp_719 },
	{ "v16@4:8i12i16i20", (superfunc)super_720, (IMP)meth_imp_720 },
	{ "v16@4:8i12{_NSRange=II}16", (superfunc)super_721, (IMP)meth_imp_721 },
	{ "v16@4:8q12@20", (superfunc)super_722, (IMP)meth_imp_722 },
	{ "v16@4:8r*12I16^v20", (superfunc)super_723, (IMP)meth_imp_723 },
	{ "v16@4:8r*12I16r^v20", (superfunc)super_724, (IMP)meth_imp_724 },
	{ "v16@4:8r*12{_NSPoint=ff}16", (superfunc)super_725, (IMP)meth_imp_725 },
	{ "v16@4:8{_NSPoint=ff}12@20", (superfunc)super_726, (IMP)meth_imp_726 },
	{ "v16@4:8{_NSPoint=ff}12i20", (superfunc)super_727, (IMP)meth_imp_727 },
	{ "v16@4:8{_NSRange=II}12@20", (superfunc)super_728, (IMP)meth_imp_728 },
	{ "v16@4:8{_NSRange=II}12r^v20", (superfunc)super_729, (IMP)meth_imp_729 },
	{ "v17@4:8@12@16@20c24", (superfunc)super_730, (IMP)meth_imp_730 },
	{ "v17@4:8@12c16c20c24", (superfunc)super_731, (IMP)meth_imp_731 },
	{ "v17@4:8@12{_NSRange=II}16c24", (superfunc)super_732, (IMP)meth_imp_732 },
	{ "v17@4:8^v12I16c20c24", (superfunc)super_733, (IMP)meth_imp_733 },
	{ "v17@4:8^v12{_NSRange=II}16c24", (superfunc)super_734, (IMP)meth_imp_734 },
	{ "v17@4:8i12c16c20c24", (superfunc)super_735, (IMP)meth_imp_735 },
	{ "v17@4:8i12i16@20c24", (superfunc)super_736, (IMP)meth_imp_736 },
	{ "v17@4:8i12i16i20c24", (superfunc)super_737, (IMP)meth_imp_737 },
	{ "v17@4:8{_NSRange=II}12^v20c24", (superfunc)super_738, (IMP)meth_imp_738 },
	{ "v17@4:8{_NSRange=II}12i20c24", (superfunc)super_739, (IMP)meth_imp_739 },
	{ "v20@4:8@12:16#20#24", (superfunc)super_740, (IMP)meth_imp_740 },
	{ "v20@4:8@12:16@20@24", (superfunc)super_741, (IMP)meth_imp_741 },
	{ "v20@4:8@12:16I20I24", (superfunc)super_742, (IMP)meth_imp_742 },
	{ "v20@4:8@12@16:20^v24", (superfunc)super_743, (IMP)meth_imp_743 },
	{ "v20@4:8@12@16@20@24", (superfunc)super_744, (IMP)meth_imp_744 },
	{ "v20@4:8@12@16@20I24", (superfunc)super_745, (IMP)meth_imp_745 },
	{ "v20@4:8@12@16@20i24", (superfunc)super_746, (IMP)meth_imp_746 },
	{ "v20@4:8@12@16I20@24", (superfunc)super_747, (IMP)meth_imp_747 },
	{ "v20@4:8@12@16i20@24", (superfunc)super_748, (IMP)meth_imp_748 },
	{ "v20@4:8@12@16i20i24", (superfunc)super_749, (IMP)meth_imp_749 },
	{ "v20@4:8@12@16l20@24", (superfunc)super_750, (IMP)meth_imp_750 },
	{ "v20@4:8@12@16{_NSRange=II}20", (superfunc)super_751, (IMP)meth_imp_751 },
	{ "v20@4:8@12I16@20*24", (superfunc)super_752, (IMP)meth_imp_752 },
	{ "v20@4:8@12I16@24", (superfunc)super_753, (IMP)meth_imp_753 },
	{ "v20@4:8@12I16I20^I24", (superfunc)super_754, (IMP)meth_imp_754 },
	{ "v20@4:8@12^{__CFPasteboard=}16i20^v24", (superfunc)super_755, (IMP)meth_imp_755 },
	{ "v20@4:8@12c16i20i24", (superfunc)super_756, (IMP)meth_imp_756 },
	{ "v20@4:8@12i16I20@24", (superfunc)super_757, (IMP)meth_imp_757 },
	{ "v20@4:8@12{_NSPoint=ff}16I24", (superfunc)super_758, (IMP)meth_imp_758 },
	{ "v20@4:8@12{_NSRange=II}16@24", (superfunc)super_759, (IMP)meth_imp_759 },
	{ "v20@4:8I12{_NSRange=II}16i24", (superfunc)super_760, (IMP)meth_imp_760 },
	{ "v20@4:8^?12^v16{_NSRange=II}20", (superfunc)super_761, (IMP)meth_imp_761 },
	{ "v20@4:8^f12^f16^f20^f24", (superfunc)super_762, (IMP)meth_imp_762 },
	{ "v20@4:8^i12^i16{_NSPoint=ff}20", (superfunc)super_763, (IMP)meth_imp_763 },
	{ "v20@4:8^v12l16l20l24", (superfunc)super_764, (IMP)meth_imp_764 },
	{ "v20@4:8^v12r*16^I20@24", (superfunc)super_765, (IMP)meth_imp_765 },
	{ "v20@4:8c12@16@20@24", (superfunc)super_766, (IMP)meth_imp_766 },
	{ "v20@4:8i12@16:20^v24", (superfunc)super_767, (IMP)meth_imp_767 },
	{ "v20@4:8{_NSPoint=ff}12{_NSPoint=ff}20", (superfunc)super_768, (IMP)meth_imp_768 },
	{ "v20@4:8{_NSPoint=ff}12{_NSRange=II}20", (superfunc)super_769, (IMP)meth_imp_769 },
	{ "v20@4:8{_NSRange=II}12@20I24", (superfunc)super_770, (IMP)meth_imp_770 },
	{ "v20@4:8{_NSRange=II}12^@20I24", (superfunc)super_771, (IMP)meth_imp_771 },
	{ "v20@4:8{_NSRange=II}12c20^{_NSRange=II}24", (superfunc)super_772, (IMP)meth_imp_772 },
	{ "v20@4:8{_NSRange=II}12i20^{_NSRange=II}24", (superfunc)super_773, (IMP)meth_imp_773 },
	{ "v20@4:8{_NSRange=II}12r*20I24", (superfunc)super_774, (IMP)meth_imp_774 },
	{ "v20@4:8{_NSRange=II}12r^S20I24", (superfunc)super_775, (IMP)meth_imp_775 },
	{ "v20@4:8{_NSRange=II}12{_NSRange=II}20", (superfunc)super_776, (IMP)meth_imp_776 },
	{ "v20@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12", (superfunc)super_777, (IMP)meth_imp_777 },
	{ "v20@4:8{_NSSize=ff}12{_NSRange=II}20", (superfunc)super_778, (IMP)meth_imp_778 },
	{ "v20@4:8{_NSSize=ff}12{_NSSize=ff}20", (superfunc)super_779, (IMP)meth_imp_779 },
	{ "v21@4:8@12@16@20@24c28", (superfunc)super_780, (IMP)meth_imp_780 },
	{ "v21@4:8@12i16c20c24c28", (superfunc)super_781, (IMP)meth_imp_781 },
	{ "v21@4:8@12i16i20i24c28", (superfunc)super_782, (IMP)meth_imp_782 },
	{ "v21@4:8i12i16c20c24c28", (superfunc)super_783, (IMP)meth_imp_783 },
	{ "v21@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28", (superfunc)super_784, (IMP)meth_imp_784 },
	{ "v24@4:8*12I16{_NSRange=II}20^{_NSRange=II}28", (superfunc)super_785, (IMP)meth_imp_785 },
	{ "v24@4:8:12@16@20I24@28", (superfunc)super_786, (IMP)meth_imp_786 },
	{ "v24@4:8@12:16@20@24I28", (superfunc)super_787, (IMP)meth_imp_787 },
	{ "v24@4:8@12:16@20@24i28", (superfunc)super_788, (IMP)meth_imp_788 },
	{ "v24@4:8@12@16@20:24^v28", (superfunc)super_789, (IMP)meth_imp_789 },
	{ "v24@4:8@12@16@20I24@28", (superfunc)super_790, (IMP)meth_imp_790 },
	{ "v24@4:8@12@16i20@28", (superfunc)super_791, (IMP)meth_imp_791 },
	{ "v24@4:8@12c16@20:24^v28", (superfunc)super_792, (IMP)meth_imp_792 },
	{ "v24@4:8@12i16@20:24^v28", (superfunc)super_793, (IMP)meth_imp_793 },
	{ "v24@4:8@12{_NSPoint=ff}16{_NSPoint=ff}24", (superfunc)super_794, (IMP)meth_imp_794 },
	{ "v24@4:8@12{_NSRange=II}16{_NSRange=II}24", (superfunc)super_795, (IMP)meth_imp_795 },
	{ "v24@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_796, (IMP)meth_imp_796 },
	{ "v24@4:8I12{_NSPoint=ff}16I24@28", (superfunc)super_797, (IMP)meth_imp_797 },
	{ "v24@4:8^I12^I16^I20{_NSRange=II}24", (superfunc)super_798, (IMP)meth_imp_798 },
	{ "v24@4:8^f12^f16^f20^f24^f28", (superfunc)super_799, (IMP)meth_imp_799 },
	{ "v24@4:8^v12^@16^@20^I24^@28", (superfunc)super_800, (IMP)meth_imp_800 },
	{ "v24@4:8^{_NSGlyphGenContext=iiiiiiiiiii@[32i][32i][32i][64i]{_NSRange=II}{_NSRange=II}ii^{_NSGlyphInsertBuffer}}12@16@20^{_NSRAStringBuffer=@IIIIII[100S]}24@28", (superfunc)super_801, (IMP)meth_imp_801 },
	{ "v24@4:8^{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_802, (IMP)meth_imp_802 },
	{ "v24@4:8c12I16r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}20r^{_NSRect={_NSPoint=ff}{_NSSize=ff}}24^{_NSRect={_NSPoint=ff}{_NSSize=ff}}28", (superfunc)super_803, (IMP)meth_imp_803 },
	{ "v24@4:8c12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_804, (IMP)meth_imp_804 },
	{ "v24@4:8i12@16:20i24i28", (superfunc)super_805, (IMP)meth_imp_805 },
	{ "v24@4:8i12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16", (superfunc)super_806, (IMP)meth_imp_806 },
	{ "v24@4:8{_NSPoint=ff}12{_NSPoint=ff}20@28", (superfunc)super_807, (IMP)meth_imp_807 },
	{ "v24@4:8{_NSRange=II}12@20{_NSRange=II}24", (superfunc)super_808, (IMP)meth_imp_808 },
	{ "v24@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28", (superfunc)super_809, (IMP)meth_imp_809 },
	{ "v24@4:8{_NSSize=ff}12^{_NSSize=ff}20^{_NSRect={_NSPoint=ff}{_NSSize=ff}}24^{_NSRect={_NSPoint=ff}{_NSSize=ff}}28", (superfunc)super_810, (IMP)meth_imp_810 },
	{ "v25@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16c32", (superfunc)super_811, (IMP)meth_imp_811 },
	{ "v25@4:8i12i16c20c24c28c32", (superfunc)super_812, (IMP)meth_imp_812 },
	{ "v25@4:8{_NSPoint=ff}12{_NSPoint=ff}20@28c32", (superfunc)super_813, (IMP)meth_imp_813 },
	{ "v25@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28c32", (superfunc)super_814, (IMP)meth_imp_814 },
	{ "v25@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28c32", (superfunc)super_815, (IMP)meth_imp_815 },
	{ "v28@4:8:12@16@20i24@32", (superfunc)super_816, (IMP)meth_imp_816 },
	{ "v28@4:8@12@16@20@24:28^v32", (superfunc)super_817, (IMP)meth_imp_817 },
	{ "v28@4:8@12@16i20@24:28^v32", (superfunc)super_818, (IMP)meth_imp_818 },
	{ "v28@4:8@12@16{_NSRect={_NSPoint=ff}{_NSSize=ff}}20", (superfunc)super_819, (IMP)meth_imp_819 },
	{ "v28@4:8@12i16{_NSRect={_NSPoint=ff}{_NSSize=ff}}20", (superfunc)super_820, (IMP)meth_imp_820 },
	{ "v28@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32", (superfunc)super_821, (IMP)meth_imp_821 },
	{ "v28@4:8@12{_NSSize=ff}16i24^i28^i32", (superfunc)super_822, (IMP)meth_imp_822 },
	{ "v28@4:8I12{_NSRange=II}16i24{_NSRange=II}28", (superfunc)super_823, (IMP)meth_imp_823 },
	{ "v28@4:8^{_PartStruct=if}12^I16{_NSRect={_NSPoint=ff}{_NSSize=ff}}20", (superfunc)super_824, (IMP)meth_imp_824 },
	{ "v28@4:8c12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32", (superfunc)super_825, (IMP)meth_imp_825 },
	{ "v28@4:8i12^{_NSGlyphGenContext=iiiiiiiiiii@[32i][32i][32i][64i]{_NSRange=II}{_NSRange=II}ii^{_NSGlyphInsertBuffer}}16@20@24^{_NSRAStringBuffer=@IIIIII[100S]}28@32", (superfunc)super_826, (IMP)meth_imp_826 },
	{ "v28@4:8{_NSAffineTransformStruct=ffffff}12", (superfunc)super_827, (IMP)meth_imp_827 },
	{ "v28@4:8{_NSPoint=ff}12{_NSPoint=ff}20{_NSPoint=ff}28", (superfunc)super_828, (IMP)meth_imp_828 },
	{ "v28@4:8{_NSRange=II}12{_NSRange=II}20i28^{_NSRange=II}32", (superfunc)super_829, (IMP)meth_imp_829 },
	{ "v28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32", (superfunc)super_830, (IMP)meth_imp_830 },
	{ "v28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28I32", (superfunc)super_831, (IMP)meth_imp_831 },
	{ "v28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28@32", (superfunc)super_832, (IMP)meth_imp_832 },
	{ "v28@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSSize=ff}28", (superfunc)super_833, (IMP)meth_imp_833 },
	{ "v32@4:8@12@16f36@24@28", (superfunc)super_834, (IMP)meth_imp_834 },
	{ "v32@4:8@12f36", (superfunc)super_835, (IMP)meth_imp_835 },
	{ "v32@4:8@12i16f36", (superfunc)super_836, (IMP)meth_imp_836 },
	{ "v32@4:8^{_NXStream=I**iilii^{stream_functions}^v}12i16f36", (superfunc)super_837, (IMP)meth_imp_837 },
	{ "v32@4:8c12f36", (superfunc)super_838, (IMP)meth_imp_838 },
	{ "v32@4:8f36", (superfunc)super_839, (IMP)meth_imp_839 },
	{ "v32@4:8f36@16", (superfunc)super_840, (IMP)meth_imp_840 },
	{ "v32@4:8f36@16@20@24", (superfunc)super_841, (IMP)meth_imp_841 },
	{ "v32@4:8i12f36", (superfunc)super_842, (IMP)meth_imp_842 },
	{ "v32@4:8i12i16f36", (superfunc)super_843, (IMP)meth_imp_843 },
	{ "v32@4:8r^f12f36", (superfunc)super_844, (IMP)meth_imp_844 },
	{ "v32@4:8r^f12i16f36", (superfunc)super_845, (IMP)meth_imp_845 },
	{ "v32@4:8{_NSPoint=ff}12f36", (superfunc)super_846, (IMP)meth_imp_846 },
	{ "v32@4:8{_NSPoint=ff}12i20f36", (superfunc)super_847, (IMP)meth_imp_847 },
	{ "v32@4:8{_NSPoint=ff}12{_NSPoint=ff}20f36", (superfunc)super_848, (IMP)meth_imp_848 },
	{ "v32@4:8{_NSPoint=ff}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}20f36", (superfunc)super_849, (IMP)meth_imp_849 },
	{ "v32@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12f36", (superfunc)super_850, (IMP)meth_imp_850 },
	{ "v36@4:8:12@16d36", (superfunc)super_851, (IMP)meth_imp_851 },
	{ "v36@4:8:12@16d36@28", (superfunc)super_852, (IMP)meth_imp_852 },
	{ "v36@4:8@12@16@20@24@28:32^v40", (superfunc)super_853, (IMP)meth_imp_853 },
	{ "v36@4:8@12@16@20@24@28@32@40", (superfunc)super_854, (IMP)meth_imp_854 },
	{ "v36@4:8@12@16@20@24@28@32c43", (superfunc)super_855, (IMP)meth_imp_855 },
	{ "v36@4:8@12I16{_NSRange=II}20i28{_NSRange=II}36", (superfunc)super_856, (IMP)meth_imp_856 },
	{ "v36@4:8@12^@16^c20^@24^@28^:32^I40", (superfunc)super_857, (IMP)meth_imp_857 },
	{ "v36@4:8@12d36", (superfunc)super_858, (IMP)meth_imp_858 },
	{ "v36@4:8@12i16d36", (superfunc)super_859, (IMP)meth_imp_859 },
	{ "v36@4:8@12{_NSPoint=ff}16f36@28i32@40", (superfunc)super_860, (IMP)meth_imp_860 },
	{ "v36@4:8@12{_NSRange=II}16I24I28^{_NSRange=II}32^I40", (superfunc)super_861, (IMP)meth_imp_861 },
	{ "v36@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32c43", (superfunc)super_862, (IMP)meth_imp_862 },
	{ "v36@4:8@12{_NSSize=ff}16@24@28i32i40", (superfunc)super_863, (IMP)meth_imp_863 },
	{ "v36@4:8^i12^i16^i20^i24^i28^i32@40", (superfunc)super_864, (IMP)meth_imp_864 },
	{ "v36@4:8c12c16c20c24@28:32^v40", (superfunc)super_865, (IMP)meth_imp_865 },
	{ "v36@4:8c12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32@40", (superfunc)super_866, (IMP)meth_imp_866 },
	{ "v36@4:8d36", (superfunc)super_867, (IMP)meth_imp_867 },
	{ "v36@4:8d36@20", (superfunc)super_868, (IMP)meth_imp_868 },
	{ "v36@4:8d36@20:24@28", (superfunc)super_869, (IMP)meth_imp_869 },
	{ "v36@4:8d36@20:24@28@32", (superfunc)super_870, (IMP)meth_imp_870 },
	{ "v36@4:8d36c20", (superfunc)super_871, (IMP)meth_imp_871 },
	{ "v36@4:8i12i16i20{_NSRect={_NSPoint=ff}{_NSSize=ff}}28", (superfunc)super_872, (IMP)meth_imp_872 },
	{ "v36@4:8{_NSPoint=ff}12d36", (superfunc)super_873, (IMP)meth_imp_873 },
	{ "v36@4:8{_NSPoint=ff}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}20i40", (superfunc)super_874, (IMP)meth_imp_874 },
	{ "v36@4:8{_NSPoint=ff}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}20i40f36", (superfunc)super_875, (IMP)meth_imp_875 },
	{ "v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32@40", (superfunc)super_876, (IMP)meth_imp_876 },
	{ "v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28I32@40", (superfunc)super_877, (IMP)meth_imp_877 },
	{ "v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28c32i40", (superfunc)super_878, (IMP)meth_imp_878 },
	{ "v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28i32i40", (superfunc)super_879, (IMP)meth_imp_879 },
	{ "v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12I28i32c43", (superfunc)super_880, (IMP)meth_imp_880 },
	{ "v36@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12c28@32c43", (superfunc)super_881, (IMP)meth_imp_881 },
	{ "v40@4:8@12f36f44c24", (superfunc)super_882, (IMP)meth_imp_882 },
	{ "v40@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16@32I40@44", (superfunc)super_883, (IMP)meth_imp_883 },
	{ "v40@4:8@12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16c32@40c47", (superfunc)super_884, (IMP)meth_imp_884 },
	{ "v40@4:8f36f44", (superfunc)super_885, (IMP)meth_imp_885 },
	{ "v40@4:8{_NSPoint=ff}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}20c43c47", (superfunc)super_886, (IMP)meth_imp_886 },
	{ "v40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32@40@44", (superfunc)super_887, (IMP)meth_imp_887 },
	{ "v40@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32", (superfunc)super_888, (IMP)meth_imp_888 },
	{ "v44@4:8@12{_NSPoint=ff}16{_NSSize=ff}24@32@40@44c51", (superfunc)super_889, (IMP)meth_imp_889 },
	{ "v44@4:8d36d44", (superfunc)super_890, (IMP)meth_imp_890 },
	{ "v44@4:8f36{_NSPoint=ff}16{_NSPoint=ff}24{_NSPoint=ff}36{_NSPoint=ff}44", (superfunc)super_891, (IMP)meth_imp_891 },
	{ "v44@4:8i12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16{_NSRect={_NSPoint=ff}{_NSSize=ff}}36", (superfunc)super_892, (IMP)meth_imp_892 },
	{ "v44@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12@28@32@40i44i48", (superfunc)super_893, (IMP)meth_imp_893 },
	{ "v44@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32@48", (superfunc)super_894, (IMP)meth_imp_894 },
	{ "v44@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32c51", (superfunc)super_895, (IMP)meth_imp_895 },
	{ "v44@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRect={_NSPoint=ff}{_NSSize=ff}}32i48f36", (superfunc)super_896, (IMP)meth_imp_896 },
	{ "v48@4:8@12@16{_NSPoint=ff}20{_NSSize=ff}28@40@44@48c55", (superfunc)super_897, (IMP)meth_imp_897 },
	{ "v48@4:8@12@16{_NSRect={_NSPoint=ff}{_NSSize=ff}}20{_NSRect={_NSPoint=ff}{_NSSize=ff}}40f36", (superfunc)super_898, (IMP)meth_imp_898 },
	{ "v48@4:8i12f36f44f52", (superfunc)super_899, (IMP)meth_imp_899 },
	{ "v48@4:8{_NSPoint=ff}12f36f44f52", (superfunc)super_900, (IMP)meth_imp_900 },
	{ "v48@4:8{_NSPoint=ff}12f36f44f52c32", (superfunc)super_901, (IMP)meth_imp_901 },
	{ "v48@4:8{_NSRect={_NSPoint=ff}{_NSSize=ff}}12{_NSRange=II}28{_NSRect={_NSPoint=ff}{_NSSize=ff}}40", (superfunc)super_902, (IMP)meth_imp_902 },
	{ "v4@4:8", (superfunc)super_903, (IMP)meth_imp_903 },
	{ "v52@4:8i12{_NSRect={_NSPoint=ff}{_NSSize=ff}}16{_NSRect={_NSPoint=ff}{_NSSize=ff}}36c55i56", (superfunc)super_904, (IMP)meth_imp_904 },
	{ "v52@4:8{_NSPoint=ff}12d36d44d52", (superfunc)super_905, (IMP)meth_imp_905 },
	{ "v5@4:8C12", (superfunc)super_906, (IMP)meth_imp_906 },
	{ "v5@4:8c12", (superfunc)super_907, (IMP)meth_imp_907 },
	{ "v6@4:8S12", (superfunc)super_908, (IMP)meth_imp_908 },
	{ "v8@4:8#12", (superfunc)super_909, (IMP)meth_imp_909 },
	{ "v8@4:8*12", (superfunc)super_910, (IMP)meth_imp_910 },
	{ "v8@4:8:12", (superfunc)super_911, (IMP)meth_imp_911 },
	{ "v8@4:8@12", (superfunc)super_912, (IMP)meth_imp_912 },
	{ "v8@4:8I12", (superfunc)super_913, (IMP)meth_imp_913 },
	{ "v8@4:8L12", (superfunc)super_914, (IMP)meth_imp_914 },
	{ "v8@4:8^*12", (superfunc)super_915, (IMP)meth_imp_915 },
	{ "v8@4:8^@12", (superfunc)super_916, (IMP)meth_imp_916 },
	{ "v8@4:8^S12", (superfunc)super_917, (IMP)meth_imp_917 },
	{ "v8@4:8^f12", (superfunc)super_918, (IMP)meth_imp_918 },
	{ "v8@4:8^v12", (superfunc)super_919, (IMP)meth_imp_919 },
	{ "v8@4:8^{?=^{_NSModalSession}c@}12", (superfunc)super_920, (IMP)meth_imp_920 },
	{ "v8@4:8^{?=ddd}12", (superfunc)super_921, (IMP)meth_imp_921 },
	{ "v8@4:8^{AEDesc=I^^{OpaqueAEDataStorageType}}12", (superfunc)super_922, (IMP)meth_imp_922 },
	{ "v8@4:8^{CGContext=}12", (superfunc)super_923, (IMP)meth_imp_923 },
	{ "v8@4:8^{FSRef=[80C]}12", (superfunc)super_924, (IMP)meth_imp_924 },
	{ "v8@4:8^{OpaqueCoreDrag=}12", (superfunc)super_925, (IMP)meth_imp_925 },
	{ "v8@4:8^{OpaqueCoreDragHandler=}12", (superfunc)super_926, (IMP)meth_imp_926 },
	{ "v8@4:8^{OpaqueIconRef=}12", (superfunc)super_927, (IMP)meth_imp_927 },
	{ "v8@4:8^{OpaqueMenuHandle=}12", (superfunc)super_928, (IMP)meth_imp_928 },
	{ "v8@4:8^{OpaquePMPageFormat=}12", (superfunc)super_929, (IMP)meth_imp_929 },
	{ "v8@4:8^{OpaquePMPrintSettings=}12", (superfunc)super_930, (IMP)meth_imp_930 },
	{ "v8@4:8^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}12", (superfunc)super_931, (IMP)meth_imp_931 },
	{ "v8@4:8^{_NSRefCountedRunArray=IIIIII[0{_NSRunArrayItem=I@}]}12", (superfunc)super_932, (IMP)meth_imp_932 },
	{ "v8@4:8^{_NSSortState=iIIII[4@]}12", (superfunc)super_933, (IMP)meth_imp_933 },
	{ "v8@4:8^{_NSZone=}12", (superfunc)super_934, (IMP)meth_imp_934 },
	{ "v8@4:8^{__CFHTTPMessage=}12", (superfunc)super_935, (IMP)meth_imp_935 },
	{ "v8@4:8^{__CFString=}12", (superfunc)super_936, (IMP)meth_imp_936 },
	{ "v8@4:8^{tiff=*^{_NXStream}sccsll{?=IIIIIISSSSSSSSSSIIIffSSffII[2S]ISSSSI^S^S^S^S[3^S]*********[2I]II^I^I[2S]^f[2S]S^f^f^f[4^S]S[2S]**I^v}{?=SSL}^i^i[10i]liillil^?^?^?^?^?^?^?^?^?^?^?^?*ii*l*llii}12", (superfunc)super_937, (IMP)meth_imp_937 },
	{ "v8@4:8i12", (superfunc)super_938, (IMP)meth_imp_938 },
	{ "v8@4:8l12", (superfunc)super_939, (IMP)meth_imp_939 },
	{ "v8@4:8r*12", (superfunc)super_940, (IMP)meth_imp_940 },
	{ "v8@4:8r^v12", (superfunc)super_941, (IMP)meth_imp_941 },
	{ "v9@4:8@12c16", (superfunc)super_942, (IMP)meth_imp_942 },
	{ "v9@4:8^{_NSModalSession=@@^{_NSModalSession}iciI^vi@@:^vi}12c16", (superfunc)super_943, (IMP)meth_imp_943 },
	{ "v9@4:8^{_NSSize=ff}12c16", (superfunc)super_944, (IMP)meth_imp_944 },
	{ "v9@4:8c12c16", (superfunc)super_945, (IMP)meth_imp_945 },
	{ "v9@4:8i12c16", (superfunc)super_946, (IMP)meth_imp_946 },
	{0, 0}
};

int ObjC_RegisterStdStubs(struct pyobjc_api* api)
{
	struct method_table* cur = method_table;

	ObjC_API = api;


	while (cur->signature) {
		if (ObjC_RegisterSignatureMapping(
				cur->signature,
				cur->call_super,
				cur->implementation) < 0) {
			return -1;
		}
		cur ++;
	}
	return 0;
}
